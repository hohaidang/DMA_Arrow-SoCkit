��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛������#O��v�,�+�v���4�ۢ��䐵I����ZG;�uwUhﺜ�i'��w�	�G�1�fV�7�ϊ�Ó���8�C4��=�҇k�M��9�Q����Ǟ�H� �a�C�����c���t/֨]�}��_il�}+�?�e�g�e�Fݰ�6S)>�>��'����Pp�÷�x�S���>���9з�9MN�V��~��a�$��5���#���;z3u��P.�s�k${�s[i��M��RԓQX��=����-�K��˄�́_��2a��愮#�����N`��r;�����4j�ֵ����=�KQ���n�r��i;�G�C���?s���|rÿd��h�eZ�ud�"?��>�ӏ��9b
^���+�k*��d�QF���ר���uQ��V?��F܌����xcVs�Ҵt
�"B�J��ʾ�U�����*�d�CȼJۉg܆���_��6�@��:M.�簨ԙ�biUۓm�j�ј_�o֩UW��?ޙG�-𥏯����s/V��̞U�L��5��g�C�ܟ_��a��ƽ�ݽ�]��H��阙#�g�����O�\�}S�6h�P���0��~���xg�Q��#�o��&m�y�+F*,�M��+r��Mb������}�$�z�ӟ�O��Q�
��زC��&����~ZZ$"����~tĆ;
�
R�-�F���0�B�')R�mfiD���F���P�� ��F�Z
Z�Ξ�:�s���~15; �󫰓��eP�V\\��"�+�N���SS����V�\�P3N�pRc?��pc��2Z2�P!�Y�X=wl�	�E��M}F!�WBdY ��%���F���;�q��L���a��s!q�7)p����!L;bp6��R��Y1���zPkV-VIe��U����#���`�t�XՎD��	_�(�e�<4?�sx���Ͻ����vl.'�|� oѣ�8�sΘށ33�
 ߭��KgC�������]/Ҋ���9Y'�\;�C��M�|r!C7�Is��P�L*�@�U�A���0����r7hm3�v�J��lM����)�����h�J��|UoB7��T�,k_�3��Ș�(S��#Ɏ�"���-��L��������7�0�EB�U]���P\?`���Be�'	�����~���(W��'e���:,����-E*�w@�2v��5��F7�xL*�N��:�sQ�@���J�-lSJ��-�eD��� �Ǒt�S$���8f�T��	늣MI��^�
�m.B�q W[�׫B2�BaMn����'�GV��d�̨P����a�[?���~�G*�����4_�^Oz�y�o>���Y�-�W�i�^]��kR8Q6�~/���B�.�� �G�����U��#t�o�N���cQ�>4O�V�3����	��q;r�'J}-��p�k0��n��s�r���m��=��k��Q�hc��s���.Q
�`�+n��ل�;�&���r���z�WR��I��i��t�KΊ��xJ���~{�u��l������	��nC��g�Q^�6���h��L�)J�#٣0sM� �K�Y.>)�P1"�C0~��[�#.�ئ8�ꖧ�d[T��/��vd�:����/1�Z5�%M��jY��ct�զ��6�:��3F����տD5˸�Μ��S����Ϲ@g��qv���(��PH,�pkC�mZȎ) b�[,��v��ay�"��d���:�J*��!َ2e�7S���W�o,�0����d�	R�r�	)�<����������j�����tu�ip����b<M��T\.�T�?w�q%�-�U�R�if��#�9���G|����h���*� 5z��Ç��Y配��t�ZXf�spi��B�\�j-g�J`���?;"�?5W��.���M��ș��v��C��]��,G�����	�z��nS�ʺ��Vg�����h������w���K��5�iҠ�ߒ�xRڒB�|��
�%M���1���`u��Ӆ����H��ս�9E�<�%�a}}j�!T�H�l�Rvר'@ //���tNP��I�SM��4������C�{Y�
bH�?�9D�`ܶ;\9��|��[hcy�o=�����9�\�!��zsQol��cY�[�k�;	��3��檛V.�k���v�C��jl/��q[�϶)���M�%V�X#�l��5Dx��c�2�k�ۃ�ې�X��O�!���hv�X���Pou��(͌�g2t"M-c�R�Y�(�C`���:�Garp��_�K��W�hg\P�E�HW۶F���?Bwߣ�㸕^��M�64�A��u�q��	������� 9������J=A���۽� ��m��v+r��7���?!��Q3$��)r���)ՅV}��P�c- 
q+�+��ASM}�t�.F��=��e�E�(/�~��׋,�te��۩T t��Ɏ���]2�,m-J���EU �'}�_4ԍ���������;�%�+���e���fd�nTc3�������qumY��� 9�9�ev�j!~�%�'ϯ��jDp����,�:1Z�<�;��9�v�l���̋���`v�A*�/C�in��^�R9�5�x�@�9�A�ȳ��� ��2���� *V?��泸EZ�t��۬ �r1<�1����0��)]�̰�]o�������;�g�/Z�}Z�����W�����<Ÿ��ͼ4xB"{Fz���P`��84G⤽-��i�-�F�)L}a��}ǧG4,��dџ�G���Z�`�W��>]б`����b7	����Ʋ��8ݐ����8qy��d�W0;PV�4�)���C6�.ln_<-�֩�01|�O�.���&�pVrL�Euf�ͨ�8�"���S�n濙D������1�α��O�D��6����Qo!���h�crt�ŭ�ۘ>]o� �P�ʙ¾��Ji�[�W>b���?
rk���)4�m�,��R_'��|�ἩW�`�06>{O�_{*ǆpY�A����?����J�B�3���7!��t��/��%��+��v���guuj$�>�oM�9{��
p�5�z�z��U��6�~I!��ψ¹��_!�k�r�z�<S���Z*DVu9Hm���7밸�WL`�#���_r�-D+PB7���ȿM�@��S9���{��
r��O����!����D#�d��:2J�֭�h<m��n�>y8M����A׸�e�&�r7(��~�/�?~�#h�Ö+G��Μ��x��z�52�;��Ш�4�)�\��K�˿� �Z ��Y�/ݗ|�S׺p]��Y�(o>y%ʋ^�WrE�E��;��̪)�Ɵ.�!7���Ե���Ȱct�4�Ve�g ���Q��a-�8
�c|�<��[Ty�%��jW�6
�~�}I���1�}�t�Z�)%���Ibޗ� ��=uU�^�#��N�C��!�dԀ�+&*<)�ϰZ2���X�1��ŉ��F��r�y:�Q+B]2�#�1C'��:뮵7)�P�*˹q��l�s�1��&�>�������@�+�!j�5r���i`�Qook���4��t�S���N�\筳i�?�fn�n���JHk�+E��v'�E����բ{����e&ѡp�>�B-���?U2����c����ՙ��6��ʲ���q(�mw����u�P!�8#l���l�U�yN����Y?G/U�m��S�&SƮ��VH\����Մ?�"ʹ̅k��2�t��*�0a�*�٨���[����юGQ�����kS��2�4$S~�Ox&�	~����v�Ο*�a?}���23���aH��Y9tK@���.<�[k5��^f�T����C �ѠWF��D�42c�$�L�������͌E@LbC+ߚ5�\F�Uљn�8��+鵶�e2F{�v�*��?,�F�Qt���#���&`s-d��is�b=1.Z<�{�y7lj�k'6V� X�����`��s�;lo�C}�;�$?�rg�28FD���>b��~�_S�}�n|����~p��ݾ���v5���>?�+���W-z�ˣ���A��'Mٹ��q��wZ�3уvd��ڴ���oE��Z�D_�0���l�͘0$5oR�t���m��9ٱ��9�Q}�L��j��C�8076�Y5$�����>������J�c�h��f��t���S4�!6΅�f#$"��!p~+6)��� �1�T���Y�=O���6�y�h�R	&V��g����B8@��77��c6�P�]���n)�/��)��y���^G��U��E��Ss����5� R���Ȇ�%�l��_\D%�t��r��1P�Q�_��e�M��C	#�c�F�J��(�{�78�2{�'א&}��U ��-\�r�#�yc��Eqt�2� ���Ο"�'ڪK��F��P	���ا�;�w���5�}2�+��4)��K�9��e��vͻ 0�������ޔ����E&��|��$"7-.4~}B,���fq���g	^�da�5��D#)�l�� ;��{�g8��F�--@>q2{Q�M��[���	O�?冸XB��I��7��n�D����~%���� V��w�j�B�'0�1x�<�B6v�7�%���~ШC����_b�6�#�%�b���ؓi�%M�cғ���nXчk �f�B?��aM�p�q���pD�Z�\W�>7�NO��Mk,o9�y�0��E���;�jB}�%t:o~�>�n�z��ä��7ށ��$�����פz�'��#�z8)�hC�'Z*�l���?����IZ��<R�T�L���4T=�^eŽ#+n�az:������ƩZ��ဍp`��I^ʛǳ���#<G9)J�{y	�/���A� �L�Y�:�'Г��	s�+d��v;�L���:OB�K�8&�t�c�~G4JR�k�ҡ��>A��J�9]GV:p8ʊ���k���΍דc���6bΈb�Byb%�h���c�,ܕJXgМ��E�~���M�T9|��n�z��Vuޗ��EX�Zů��*6��ٯblEu���s�:\�SW�����܋ػ��&T��x�-9H��<�3��\���@AJ>����$���+�7`O�$�!��K���*���d��R���X>}k���O!��L�.窽����h���Ka7f���X���[o�f,h���D��5�<��ܠ�(!��6[q�8��x����_�}�ؓ���Y_��*)����@�a����1}���/q��Ab:'�s������f��5
��R�Z�����V�V�8�@+������%�:�O^HM*P)�/� �G��d1�����j'BNo���=6���BX"`i����.5+������wFV��Bx|��tM�=a���Ǌ�%e�CJW�	��`'��dW�|4#�p��
E'�3c�)�s�G��©r6�S�L޴o���
�ϖ4��;x�eb���6�*�K �P�-�3nXC15X�C7:�ǳ�	�eLƿM�|��ExX���R����a�7�
Jk[s3�Kv�ٺ��D~��~���2(1F1s�`��+��G�NnS�i�$��h#H\0�j�?�p�ou�宄0���i���Ą����l��7X�V#�C!cX���S��N2�5EC��gw⵴������M;��#��óKh�� ��x=���S
�N�o�١�[�.}/��F�(�-�d�W6<_�%�}$"
K�OT�}�z���n��@s;�ĚC7���ZUk
~�*��:,,/n�����es!o�b�����L#[@j�Z�W��3���T �'!���B�_fMe�~5y���!����,��/�p�[�
��L�F-2�Yf��������@Zُ"q������w~�[���Q*A5�����v�>��� �:s$/���+�2u��Z�W����Eb&��a2T�&�8�F�త`��7Z�N�9���������W�<@N�
z�����aI\�Z��Y~����_Ym�������~;��� =j�΍�j�ĳ|zQ@y�>%�m��?нg|��"a.��SMl�3��w<���l ?� Πv^h{����o�ٕ/��aC@��26�����Ϝ)%�D��\BW9Z�Cۺ�⼙[��faJ�F ���B��>\o�"�]�w��s%��dxv�hbE{�c�G)�����2G�ږG����l�N?�VL[����_j/��QL��U�35��u�뿲�l*���G/��L+J����DY�ˑ�5Y��_����"��St����U+qLC�}n�ܓE.qMK��<�N���
@���-�N��m��pݿ�N���^��n'�#�m�W��EE���8?�a�y�ŀ��I����:gjh�H�"������z2ǥEFE=�Ԇ������*,,��;p�x	�r����$9��ax+��C�#����JL�:��P��;�6{���ſC`^*Su���
܂�tTi�@)�zf���h�;�����3���"FȒ� �uW�ǁ�O�I���%����-��0V e�i�V�4�L����zx&O��Gk��-��K�ޣ�\�S3� +)�����$@W��t�1��� �ټS���-��"�:�0kq�9<S�o)I���l�.2g��m�Kw�%#�� �����M������B��E���k���f��C�S<�Q�����I!_�A�S{d�!R6�s���x�n��jBI�������z���ao�yf���Z�|�@+�-i�w�Nn����g�f:���E��\��r��Ï`eP�;�Y�)��i�>�Gd���� :ܞH�ɴҶo�(����d����l���R��U�Qlډ5��o�QX�v$�5��EX�C��7�+vHS+`�,� ��A3�q�Hm�:j�Gg�,�b�a�Jͼ�� ��I`�ME-�f����z�R�z�9�]��ڵ���1P��p���J��FD�S���B	�Ȃ#�wO��#������2Ғ<q ܪT`�i%���q�B�n�Z� \��������R��|�z�vf�(���:+�+�7�%{�~@�Q���ug������8|�q���I���� <�E�ԇ9�j~f5�Xz$H�5��[M�Y��ʞ�3��]�n�,��%���ʱMD��`�����O���*�ƓU��n�P��d�Y���p޲�3�/���l�V�2�]���^	\�mN�0�|	�]��L���q�[�>�0M��\犞BM��3{XƘT\�e�3��QQA�J��,�6��e���2��  �8���i@�T#+:C�ޱ��|}TcR�{��E��%sk�5�ED���fZud���~���=������Z�
p<6W����On����(&ԩ��	>���q����D*�@��[d�_���!���I�O��ɹ�ڪM�?�#�WV_�1�="�s�&K�+�ϋ:��	5���Rnl1twI1�r*Y�����o���U��"�T1��OG�-L������*��2V���-�b�1�"��������n@t�Q(�~��+8ˀ��w���&���A�#r&�F!+ѿ�OY�����Һ)��\^,T��}"A~������My>8_b�quwe<�sn9�8�q�*���I[y�,���_r>e7�����n���*P��H�Yz��ދ)U&o1�S7P�)��2�n����& Y����8X,�ǃ�*F��>0߮Z���y\�QtGB�7��$��͡��͸"!��iN�%��G Mu�mA�*��z:���:�D3�-�G�gĀ��:��𪭛��?����m��h���g��	�ePyM�j
"�g��/ � yy:�������:s�* ���`��8ɮ��P�[���)�J�Wuгd�ҸQ�c��t�KjZ�[� ���Χ�+�w �f���d�����c<wY��m~���<�q�&��o.j�]�A|[�sȍ�2�	 ޵���!���kDR`�I-�:����#���q�l���K��&J(t�#�(��{��_��)��WL\E��m��;�I��l1�vb�
�(p+�X��9�����JN�>	�VqPx0�KS�m/�sr��|�y��0���@6M(�A&ц[���I�c�Y��hQp�n�nD���������e��d?�B������0q&������_�>�xs��f�"�ħ�1�[��Y��~�8=������6]�N�c��U�?���+�m���H����e~�7�Y��Ġ��Z�F�y�3����̖���[��B5�$.�*PPd�O�UZ�U��-��΍��)�\� ���,^I�����5A�<��� ��p����?ȩx��?e���R ����%dpHv����9B�����N���!�B-L/S�XE҅��JIe/y������?���ő:��܏;�SLc>��ѓ�3�@uX͑�զ� t���O�$�Ag�BC`x�r)�i��*�����	�b8�j�}�r��<-b��&��*GU*,�q?����8������֜B D*����Ѐ/�s����-�Y}�n(� ���#	3�mk����!_����߱7����Y��4e�OHEC��.R�jmjF���]�_�Md���]�A�����Y��BV璋4Y8�N�q�W���&:§h>~h ���׋0	�G������9�R�5�rQV Q�� ��Q�+�	��𞇴���W�%�{�g�7�aȒ5�
_�;l�t��@;�n
���WD�qJ{�܁�}Y�Ss3��a �$sΠ��.�t��c��~y�0LY�Z�S��gn�T�l�e4�V��?��2&�Bb�������rXpM+[P[A�Z[0�䅠/~�H�>�LX���{6߁�|��A�s�u;����ķ�B�*��`4=���W}m�;(���y�е���H����{^'�W�Agc[����r�3�ȑ�	t� G��Ϗ��3�Vm-��W򨽅��"8�����e>�1�c����.���a!C$$�s�(��Pm]A�L}= � �B;Al�#��K�+� �b�{Qzm��:���H���رk�^�/����LP�e�_¢ԭ!�Cfi2cOx>�'��W�K�L�U��)�~u'�K��/����WW�CB�,�ޓu��%,��|� gXY�c���A�K��yV���8�6N&R�u�S^l�q(��8;��{-cܼ˾�5��N]TkLS�:�
e5�G.Kja� 5Ь#��av��G�qS�Fj㫏�C�`��xY;re�a��QH7۴�5�l�B]=O������(<�jnh�H{ӯ��Q��VDc��7uM�c�\{��n�P�"��9,�o��#A&�Z�'M�o�_�_�%d�s�,��j+�8��*���%�4g!YR3��^��B^G���e�d�3�� �a%�#E���v:�`%=?��o�0��{��B��nn��<���H̒nm�xY~�����Ef9E����������D��"��Vrn�v6��_2���T6�q,���]-ӛ8_j>��J���'�?���2a@������3n���s��d�{��\2L-�[n�(J�n���	N���f�p��<~�"�x=I����@�0�xXT5��Я/e�������ך5wy|���~�j��h����7A�CNQQ �~��LpR���I]��ftЀ�s~��:��m,[T��^kL�$rD��U D+R� �]L�lq�&�Jm,AM�(Qo:�ݷ!���,�o�2�Q�%���R�g��aU�dp��n)~�q��T8���2�aW�"<Я�uyV����Uc���������(��
B�
0O�l�@M��
�Zs,z��f� Z(��r�7��������A����7J�w�wԘ��C��<z"��lWO���?Գ���C����2��ۅ�!x�9=4������?P%�h�<|��|�d������vR÷FV)X�� p���sȜw��35������ע�������P��kx?<��+���2�\Ik?�g���8*_����	�S=�ǥ,����֌�����x�a`S0ƈ)������0���"v����H���c��Րnf2j��R���sA����V���W:9rG[5�ZNB��V3�J�V+�,�������U���ʽ\:�_�(�~~L�D�ԛ�yj���iB�`3�T�J� 7�Q)?H��T��@���fA���f�I�p��f�zj~�<��ҕ�p�d+c�?++p(F"b@f�G ��Bi1e�);�?�����?M���e�l7�o�&��@�Ɂ��T%���e���4Y�U&������~Ѫ�nf�Ǳ��1ݓ*=^�� �P�FL�ιߞ'�-�;�b����,G�!)Kw8��	�/t�Em��_b�I�-#��S����2���jK5�Ƴ�|vR�&���
�P���1''��8��K�#ѱ�Bm�6���.Y�A\���3�NAS7�աT�/n��z����n�ׁM�|<nx!�p�h|h�U9
��"��q����Y��J�Ҝ�r�$�S�B F{�`^#N�}P{��"Urk�i��旡�Ѕ�����՞��A��<z�W-��>ci��OBe{�,��>�Gz[�{I@;ev/P�Az 7�`���`ݜ�R�h4�l��S^�h�f���&"@����� P�)��Fs��9��<��0���4,����-��,���!�!��Y)n�[�z=��,#t�5n�t�˼��sg�%VR��8i@pcǐ�/�[}G@�d=�[@U�Fd4P*+�MAK��\��o�g0;2?ס��=� 5�D�c��;9Y�ς-����&�%�P%uVǛ�����y�eÓG
(��� �\:{�U�E��[�r��Ǣ��H�o}�#w<#��u����ӝ����x�]U�);T�Qʊ��Y�48g/Gz����s�|���v��\@Hl��f��M6Ï0����r�>��(yB^��
MC���܀9TU��H���J����l�S��N��d �U�ߺ���z�ᣄT*^V� �/"��ϔʾJFđ�'���Z���ST��������7q���(5�[�WWW1}K)t��QH�x�jXs�?://|����հ՗ ��E�Tz�����P4���p��,������~S��rr�㪼��zi��� ��x���姩��kz��p�}�:�?��M[�RE}��"s��\��o�okd1�,4@���^���C��B&��9Y��:��*k=�P�x�w�ŋ�]9�H7vn��~緸�iz�p����e�Kh2���2-ӏU�������h�;ٰ�c9iL��g�7̂y�F�\�iꗸ��{n�g1��c	�R'�<(?���l�3��W�/L�
! �!��������b�M�M��w���������<{x��yM��jhEfrH���J+����v@�6��`0��|+�Ǯ^P,U�xn�L��αfs�N�Gu�!�[B���V����EC���<]��Ev)YΚ-��>��Im:9�!8�i��l�f(2�V�X���1��کc!/1�VS�Z_mc.JvP�A�0�x�5��h��>��41���T��:n���O��p��G�q`�mѐ{� ϓ��t��MIXC5��J1��+jt(ϡ���]c�ǈL�J{)�إ��9	������B����R����E6
���2�~�fS�>vk� ��m����l���hxM�� ���[�~w'>v
 H�\ KMz[��e�g�c6g*v_\5�z��=_�?��cϭ��!���b��L�o����Uf��p�J�:�
�qm,p�^�#��H?����D�7�����A�BnS�?�������K���D�pB�[��6ޠQFY|����S��3��B�;��C�3w�Z3|�Ե#��<;��������wʊ�R�SF������j��AɊ2��<}���xh;��G0al@v�\F�.0��TrG�\�cK_y�Q�[����&�Y>_��<6��Q�z]��OS/�L�y�3�D��uO%c�ET�wjKI��=�� �Sz����}���(����d��Y������+�^�f\?m��oݺ�X@�ߤ�SQD$�g�a'"2bH���%kxEy�h^�kY�]1n~�Cb�SX	���%�S�ɕsUH.�Y�h�p���r�Z�j��rs,qt���I;d����_��;e��o�����X���	�B�/v�x֒�[;�f�u����V��YI`�L�V�:�׋�C$�]�~x�b��p�)��T�x�O��#{�l�Σb:�y�5Q�b��5d�o�0v�U΀x��ȍa
 [���md�B9���>Q���w�jY�m���3��yh�y�c����2 �To}��kE�8c+_�pۮ�q&�C��xR��<��t��iA��'���	�a�{q�T8�AA������Z����xR��#�ʜ>��~0�:�v�.�&A���S���uĂ*��w�Xdk���C}����+�|��"�6����,9�VQcM_Τ���M��Y<rՌ��J�PZ|0By�a���[  �%��Hk��[IB����B�i1�`\��bN8�[��!�Cl:%�Ҽ���kd.j�E*�{C<�;���)���؏dxdگ��p���gl�[�YG�ژ�)��?�����j/E������PUth�v�nY�*^}�?�Ĭ= ������iK�+��q!��D1�+��ðy��]�c�M.?[Q��cv�(��l�=��u���,O����h����v(/����ȓ��\!�.-$m}�^J�]PL\;�͜= E҆�>�6�La[6:��!��C�z��Ig'�����:��ݺ�M|�HG0��O�e��� Y)E|qb2�ou^�o��դ��]�a�Mل����@%�}n�}�(V���X4�7*B��w�U�?��������~�H� 8ֵ9?�{˅w��ɘ�B�T�Kw��2qi��Ǌ�C���(�������J�bW!�.�g������d&_��d%�d��J�F`sw�X����x�R��*r����G���o�[��q֞0���JA�-���DQr��-���&C�,�u!0�[� ��r�0g��`7�`���E�3�,@Lk�����G~$�jv�/�G7�#�J�:t�7����Yi��i<�+�-Nk����clPL�<[���Ur!�7`H��r��iK�:"ڏAC��ʿ�i��-n��n�4�Z_2�Ȇbb�lƂF9�3��۝�'G�%,D����-Z��5������ȩV���o����-!'�XI�R����A��|
���RCG-�{?��p<%�vif��b�n�]�5u�İBx������S�0�.�b�����8�߀�����������������r�5�,X���&�ű�>�F����^D_�P?�Az#jp�ؖ����y��6bU���5>cP�O�$8̴�g���ۿ& ������E��x�z�>TVI��z�+[�զ�E���D�|Bҽ��f�i͞\ �7J�W�x}zy�E����L���[\0�{9��cc�2kk�p*������/���P���F�02$ڽ���a@���@�	Y\1��/���E-�>��풀t\ j�t��m!>3�Wp� i���^�-�&��ê������ޅ��"~|��O�
�TJ�}tѡ�������*�dDAh����zb�0�V+Ѩ	**X\����mE��DN#���S�%�cζ�QY�	�{�D�J�k�%6sՒ��o5��-�H�.�_��l�Wѣ�$��0U����P���*FE��WPx��dH=���#u���X�RgO�X�gױ؍�0�x�{\��ֿ E���qz[����*�DB�+��=�O%c��w�]�앭:����/���O�j�	..��\�'İ8d'�ݡ�����G`A���3�q>s�la�ۀa,����<�
'�Y?I����\�v�~B7�����c���
;����X�HC�6�uk�D��X:�.A��186�XD}ڱ��4X��K3�+�D2�X8��`����2��!9�2�lo���C��CͷiN�?%<�\;II��AR��E�
d2�@�[���	r�^͈�r}��~"7V{0JB�5�8��^MIMPB��;�tV�E�N)��c��zW+��!/1���
���EȘ��i�j��qi��N))��3�FV�f�� ]?�m�~X���<1���#}���<�1g-XTD��s!� �n�p�uf�p(���6�wED��"���d�f�O권����Ƹ�'��R�T���l$t��H����π�D���"�ɸx�5���2��Yl�<y�ϐ��_��!�r�3��qx���lR���c��|�:�ߏ�;��.$�<E�h����7��OZ���I��u�T�Xs�f��;�v��U��3�r���H3շ��ހm��~5���ݹ�J/D�~:CG�R�F�Ҫ(Y��vYH�7��g6dL�n~�Y���:xZs�N��}�B�d~_�аG,�m�pOE�ҡ�|��3;i"u�6J�x���[�4�l���^�S?�a�*Xe���g�ne���)e��%�����9����mO�юǉ�+7�[��F!�G'��*	�o�l�����i�F�\(�t�EknpS��L7>��n�]]��<�<���\<��oF�sq���#F%�I�O=���G5��0�@,j�*	�+�����t��W"#`�'��.��[,:A��̕rx���B�V��O��T`�q�+�
J�Ԛ��b�8�Iè�
�����E�.�w�S
b���<�?�$ًi��2��=����6�#o���U:Њ��n�Z����n�Ճ.�+��1e���קO2L��y����/dII�Qk��UP�_�{x����֑օ<-Q-�E`�������.Y�W��y��������ؕ��5t��S����T" x����/��;�<�IA�^�p����T���I12��>��j�������o�"�x㪌vHm�� �������w5}@�B9��ylH����`C�_��"�G�L�*Y�R[D|ǌ��-��a��7��D�:V����7r�K����R��zX&�sR�͇�����Y�Ph̚l�3��lR|�š���F�������}�ET| G�P�DE������LkOu�z W��K�O'G�4���B�����j̐�R�ީ���Q"��-�{U�^Tvq!v��.�`��BC�[�s9�
��vš	�-m2���JL��ܯ�v��C�����k�S��Ец\���q��kT&A��]MMH
�V���D�+�5� �}B��2MG��#����ȁ���y�Yx �b��)[?{o4��d?6>���PV�cR�99B�>p��A8	D�s��u�I]6��/��ǽAOd��%'�<(��7��!�9��V���t��y�D�����
q���#�Vb�Īzl�G� Y-)<?��϶*ea˻2�����3X�ޥ{�W���8@�Be�� �iÙ�֢�W��
C~B��se���\�ì��C:)��8�Z����~LO
2%��Xq����4!��������[o��g��A�Ckk�1z�j��q$O"0f�%Ne��{V�������N��я�j�˷�ǝ����JWձ��9Ly��#7�L+�3Ƶ�S�r�2Lߺ��+d7�^�����7��y��خ)��eY�W���Q�ײ�޵ B�\3U�'d��	�U�(��zCNj��n7���N�z ��\�B��9������w^g��R��{�?߶QR�ל�RV������Էc��4�	�<�N���7?��[�<b�b��/���Wct^W���q� ����Rmhn������>�!��v�x��V+�f�n�f�q��B6�@��XN^Shb��Q�h9D�i�[6�4D��P�3� �s�>.ǎ�B�UZ�ԇ62��jh$����
��V������ȶ*R�$��}ts�bUmj"3�w��}���k�*X(�}�R;�YO9�%�/>�8��>�E�\�����=�]�3�ԁ%��ab���Y'�f̷�g�1p�<uz_IuhnY,�)O�G!dE᪐�iN��#�;�-�Ą���j�2�|B��LpL��Դ�f��ԉn����l|7_H+S���t��nJ�탑��acI�35H�0s~���Ͼ�G&M:e8��I_t9�Q����bH��I�	�n�{�Jϲ���7����ai�7?�� �w���:cL�Z�����L���f'������3��K����P���.��}��*{{v��=��3!�˒h��to�6���lEAs1�-z�����W>V���d	�EYRR[���:}�4L3	_���z+�[��&�9̩wh���o���s����<��
F��
�c|��x��ʚ��z]ո���L��1?�a2ȫort��%S���G]�$����W��v�J��(�T�}�4y��!)s�I�st����\�I���
��0�ϊSȝ���Ŏ���h��b��Zr�08bߗ@�.ȯw�U���ܒvˡ��%�\�{�F	�u��;�P���?��𲞏��A��
3�Ew��O�e�$��ȏMtQ,?������\�ii��!�9�-g���%��?c��'8���U#�xY//�QqY�����ŢT�U�s��/ّ��0S�}�;���ie��DM"��T��l{?h�����"w��Gmʧ�Z�m����"�Y�>���H�V�|퉵�p��d��E,ȩ�F�^n>O0��2LS�'7���`� ���k"��/���	��9�u5	�?1�Y/Ws׬��$����E~B�0זm<�o�^}��$�%B�o�dt��%�h��������,q����6Y	�'���J�h�n3-hБ�lz�ȟ�E��ѰP��JOS��ˀ@�ԛ︥���z�$̴� ��U�.�ԡ���V���0����_��!|�z�?��@),�����
�x�/����	t�����wZ���A����DZ���I8��泃Y.b�Qp�["�ԏ�u�(�!�aJ`ƌa�f�>�2�'�V��7�9^e�a�8K�5�V����-
M�K9�W�Z��A)��*�Sj��(��E� DC�~�1õx��d�G}��쇢�6ӕ�R��%ڨ�&9o��j""��Z���ۊ~$K��tp�ζ�g��`�-�x�fݥB󓏟7�Mݑ� ��I�.�hT��Ǫ��%'�|K�P��鵪M��:'J�!�iy�Z#����]P�{J�������G�ѣ���GO�Ua�m�����$n��v	��D%��(��F?qC]��U�f����i6�B:�M�ݓKJG\;�g`����!\\M�	.GS�k�����C�'��ČO��!���L�����㜑:���o!����}���������9 !Q
i�G6�r�c<X��Q1w����i��!L�É�8� ߳���T	��N�_�;���;h	H D�
�n^�i�k��������U苧�ˀޅD`�pH��+��[A�j]! qU]��:�?$@w�U}}{N*A���Z����`=h=kX8���SծB�p���m���d���k+�~��c��"o�5�b_^��؛�u���6� �a���ڃ�A�	��
����#,g��۬S_��Eu�9�E�}�=�#g�@���E��"��|f1�G.�+g�*լ.���]Sze��"��g��:`����h��BC�-����%����M�bP�Dl���7tT�2ap��β�����Lw�8K��S��q�[����*/���6�"L��
\��,Ǽ��4#i��Σ��A��-10y�20W3�.�'�'^��O�+Q�_:�#�BNd�S�!/��cv�4�J�[��s��/�&��so<`�I�.�?�t��������pm�8B�@ea�6��,�Gy�d�����Xe� �о��Cxg��r$QWB��-�A��5�,S����P����~�r��Pc0@�p�<˙���{�4�^C�(#:�U�B���,�Y�^Y�<F����
�#GN|�sK`ߠR�$N`�,�$;�R���Z��1��ӕ�d2���+����_N�$Ħ�S>.��У�f�3�:qQ���������!��Q����
t��#,�� �|)������V���i�v��\�an<������}�sI��u��M�	!jc�s��[16�q�F�����7,ٻmeP'�#�ow���~��	�@�<.����E���1p�L�� ��gy�?�?�!���l/W��ˤ��]?�2�jtN��_/ŵ��`mg�$D� ���`����l�C�H�i�mx�:�)�{n�-�ƶj~�UƮ��Ȫ��=~C������nC�
Hl?�&�m�Z�s��9?��_�gs�#���B��T�ŉ���<���[����]�:8�9��	^֮��Q~�`2��P���GP�"�m�<���mj◲�����q�\yɠ�xF]'HS��Yq����a�z�Բȗ���^H[��@�%ф]��jce��{c���i�п���A$<ǆUB90�����B�^sS�C��i1\�,����A�Y��^��e**Ē�&����G��@�ƈ~�.�7�����A��
Y�kŭ�l֗��T'G'�������ͻ�"H��2��:P��Xy������C�ƪ��� �F�U��Z�j�1�r�ks�{!�=�q�t�Jե��*�Tܨ��3:	��</U:�CR�F�ߙ���o�KŃ6�)a9F��ɃH��U#����,j���N��)֪�eXG�L��{�vZ��~#\:��AQ����z4�B�@1y��! h�3 �D�uͮΙ����͏�V�k��
���t\il���/H��A�i�٫�[SV��N�z��J�~��ZҚ(��H}G��IzT��kme���w�By�u|s�������d��+���f�v��)��#-�9��1>p�/�NLz_�O� "�@ �w:��ȯS5;��c�7#L���D�O�g
Mّ��P&����Vw�x���I7>�si��1�~��>[r`h~������-w���y�ip�ײ?�l��%򓔧Ft�È���.'��D����V�v�f�8��^J����B�(�6��*�en�@��Ɍ4_U�Ic7���.�u��6�H��/�;�������.H�J��/+^3W`P[�6�+R��ʽ�E�+y��-�A�b`����3�NbcL�cz%�o�q���J�g)�y*ҁ:fj��+�' z��@C���@��u9wEhsӷm�%����d� ~�UW�j�`AY���XHj�;�ո�`4��:E�I-�m��`�4p|�T.|�r�?�M��"���5�Xb��J�9��Y�/c+D��dļ�h�@b"��[��˙�{�l�ˋ���L��5AAM	<�o C����T%�����-Kl+�X��.���A�<�y���2���\�%	a���f�r8l�q� �߃	�0�1%t�r|S�v@/V��Ț+�e�v;JY�����B{.»{⬏/��q99��h�Is�i����q�՝���)TE�D3�~<ˤx#:�-�a�u��D]�rմ����	���=���m�� ���H
O�N{[Pk���c��3�,J1cyyR�y��nm�ss�s�=p{
����G�k�����
��.�����Ʉ��Y@�f��Q�b�}hE�f��GuQU��&�Q�e�4�|a�V�Tt(�R������S��v����2�GOmϝ�|�M�:en�Qs������ !�{0�"U@��x$�Q,$�U���L=�,9�0Ds�T����a2&l,��ja4�ZTd��S��\�?��� 
��Κ�ZYֽ6�K���N�w�[
��,z�֭S���ߖX>��b���E0߃��7xK˯m�P���u�VJ|����t����. ���g�����i�0C#>lF'�K�Qj����P��3�a��CT�)���*�� ��r6���>��{h�[��3ٛ hr��1�cƣd�c�y"Q��gvsd���9�#��6�5���иfQ��`e�h�aP.�Z��`�K=�����R{쮊S RD�
m��Z5���+���m�����Oq$��Km�*��MD�����j�v�0q���Ƴ#��p�]�#r����Hy�(��Z|R�;}`~�7�j771�N�����]T�؊qL#T+��y��[����Ť�2>�bZ�w�����1�l�5��X=�\󡂻�lB� ��*=��%�����8�|�_,+=�fnc��{���=5�0$�Z��AgR��B&���OQ�%��۶ 	"��\!FF��D%�0��l���x�^J�i{6]�!�RU"a�C�)�Ply�-�"�lB� Ȱ�F�6�����0U�Ƌ��$��s�F�}ke{+��wѿ�q�Kb�~ ����p"�Z$*Vs�i%�����S��H�f=V?��t��^P`{�/���4Un#�$`B�9`�kأ�ԟP��O����%i�e,w�Ɇ��O�O�j�_F����z�Wc2]E@�E�[
�ɻ����*��j�
�!
'+�}�3t]��4�d����K��:�{�t$Sy%MC���������9��lB������Բ4)�܌'�@��}��W�q�"���L�]����@��`��n��Y-D*}!Jn+�D�w/��x`0�x�A����`-�&�-��	|e_�J]|�醦B� �L8 4qp������+�El�u�w���N�9N�,���%�|�55E����6��=�D�.�n5�U5٬-�J���az�d�,�P���5��v���M�#A&K�4��ו��h`�C���ޗ�(_�}��{	��M��#����PP��7}�l4�����	�X9��젧�{��̪�8xaT5���<�dF�zɴ��đ!Jv�g��xpA�%�����"����*�jB�bD�3����e��Q�`R��%Lz"�?{��	��A�(۟7orcqXepŸ�4d�S�#��Lx9JǸ����I��X��oګ�!�P�JР�F�2��(�2��̳=�A���ST�	%�3��z��o%E��B��a�m
��DI3ή*�h?���{!�93蒼a2�pR瓈g��T�(�������w\���d}���`X�~.��& ��/�t�B	^�Z�/�PR�>~�C�ʊ�IP��r7����8�*l[l��v����:Q����S��2�B��j��U6�Wzv��_�A�e��7!�$��W�Ό���̖��:�O-�A'���:��%ݣ���0:�o\m ���+���s�a5����|Gv�{������D��ߖ��P��F�;]�]�G3&׊������f&��ʞ�?�r�vP������c�������ꇬnHȌw"De�������m���4���ٓ��絞ԋ�F\�HX.��g�� H;�T0Б�yq��C�Jk�$ь4R�ѡ���+�fO[�č��6�����2å#	X�ާE���5#B=�0daT7t���yu �c�n+��X�W�]-�PJ{������AD�R>�qH��$��8�h�`�hn7?!���S&��܄؂�Hh�ۓ�9��s�>{�״���/�������=�Ō�����s���o2d\׍q�� �K�lȮ����~���eG5NÔ��k���zQ��Q���G��AЪ��1~�TE�x����?��&e!�
�ND���޶B��+ԈZR�P�Ne�he&�ϩ���A ��@�W�C^Ϭk���q��?�^��������H�f�4��|�,e)=[�|���A��r:~�!�S"��	|��̾�Gy��Nj^K��}�K�Qrӄ��E��i�!��1O�̕���@�u7h&���Q�ӔiG�_�X��� -F�1����F1X�pb9�>�v�x���R��ٍ������]��3Z��f�@����_�#��3z'Ml�)ւ|��{Yp*�<�G�|�{wp��IVL���4�����ٴ&��U�.#w�*7�	 3h�/�Z�0�ɐ�t
�Ka�N(F쮽��!��%����6vE���^3P�wK�Ɓ��R/O�}�U��t%S�Z��C�S����os��?]O3�S���S�iN��YsJ��g����0(H&B�lY>~�f!���z��-�[�I/i��Q&�U���ha����<m�U'�◭!;2�]�U'i��I�>dei���U�o��AY�'}�<A�p�%��kH�^"W�4��q&�a�/<l�vX���`ur��cF�V�ؿis�>C�g�����80~�!1��!���7�#�3Ԯsd:3����� x����0��:{br�<�aL� ^�y�p4F-&vF4�i�NSx7�?XV8A9��4�aF��>d-!�}�"�4���㋔р��m�^�41;�A�9�T���l��h��$~��褣���az�$�>���M}5��}K F?��yɠrJ��C�)���E�u�3 �%�eW[��\���p�M��� ��e{�� ��xf,o�{�:��+�Sm����<i�ad?���d6f�����KԆ%�R��H�r�����'��,΃H�a!� �g+<�?ih�sCn {t<�O�����1;c�|��[Z�} ��i���Y5�J��`��:���J:�.�B+/P�dZ��	(���	� �_.���EM֓5*a��� I���9��}���T�;�������W-ָ4�횿2��� G9��b��,����C�5�{�k��K�(�����7�R�5��lԡ�c�2��T����@_����+�V��i�b�U�*J����X���"��������8�U|"�K4M��1P/6i��n'�o䆸R\�z���컏�24�w�Rݣ��߷D��C�O9�f���h��,gPLvA;7����Hf& ��τ0e!-�"��#�}��ȭ������F9�w����O�K�K�k:�i��p.[:UT,��o�#!QW:�M(Fƶ�,�ѿ?��H+ǃ6lb7��:�P��ڄ� xP�X�Z�At��uC�I�u��έ��E���s��6X���!C��������!�A�%���������u����I	�Ď8�E�����K�r����[:i4��dj�5��{<&��,���$w���`�����m	;�z�cS;�o@/^�t��;tCw���?Lg��Z�W�X����D�_��o�CI��֫�m��C�KsM�:��W�����3�^;�9e>����d�W�k{=��L\�:(I�Ml�CWzm(Y���$B<�J�M�ݤ%�v��s*�)E�,̘Q֥Q�'��5
���(��W��Yr�p$�%�%:��2���[��+f֒(���n{�j��u��1 ���v16z�L��D���f�co�m���ڎ�¦����c6R	O����c͉�Q2����<�W2��<��[�۰h~�~FZ}�G+����T-�����ƶ���r0��%b!��;�B���TG��7Q!�夑M�gs}�L�!��:�CWc�B���d����n*�����l�5gpo�(H�����,�V�dm��6 ��G���e|i�:P�H������]�( 9^:j�,��,�[�M����: r7}�[���3�<�*υ"�)��JvT[�DBig�ھ8X2�Pi�
�4r�Q��v��K������,[7��L�g^����1�V��]S� ���*�| 7-��墴y�%���J�>��u�$�&���s��J�m�08w̪f���_:�a�D���Ĭ�0�bVL��V�jq�F԰����'A��m;��|�R�A�����n�5]���>0�#�L�x�a�"�ň�����W3&&�jĄ���:���?���7���9޻!Q0�8�So���5x�s}��Kqo��m}�7D$&E�.ڤK�*Xg�WkAߍ:��gw!����(K�-�
uN��M�	tX6)����2 �C�G� qa�Y)�kMn�*�#Bw��� ^I*-��okH��2 �qD���c�
��$���`�g]=�l��#���^���f5�b<tUw�V��ئѳ��Ah�wl�ƤG�.��ڠ�T����(3-ӟ�hy���HV����:�`7o/lW_/ �K	��8$�1UF���S�l��U��Vo(U[�(�Λ����i|Y��m�↷���U��s�WY��K�+�`R�+٬7�z���y��v,W��J(����$��l��	2�ݙ�a,��됼L(�>�Y��8"���;-����;�B�B�zM�Z:f�L��?!���t�H�!m��}tp?�!݀�#L^*�o�>�˜� )�VZ힖8��R�,vחyb����ti002����xO�KE-�������2|
,bn���G�&�
�/��=IY|/���}�d����H�M���M�3�6nuW���Ŗ-��3hXOe�C �e»[?�!�	�v+���"T��n�8�?�w4��u�6��.\���_qM�̃F�r��'�s�m(��f�b���;���R�?�W2Ks��$�]K��!*�-(9��l̞����]���[tP�Q	�x��.&�6������+�#*ekj���P��gk)A��Y)�$`'(�1#�~�d��ܡj �2�#��(�|�4�N�Q�=ςz�Ӈ�Vx;Of�[��0%��%��m(�]��i�J�pְ!��mQ������-�o��qu�V���
����w��������i�ֲg6����ö����\GYy��˓y/.�P�R��.��W�5�:�Kd���e�_L����p ����a�o�ͻ�z�ձb~��.C쟓�SJa�db��0z�uyD�Y�X�4�D��"�y�&��/�^�/�� (l�{G�"����{l��~��D�M�oGk�Ȋi�j�VJ_�{��l\�H�׺��'�N� _�>e�#�5�8�¹��6Z��������������PH�]W;7Bd+@��ڮo)J\��~Ǆ;� s��Ìr����=@8J ߊT���/s7�d���ʢxn��
���Z��O���7��R��W"� ���%d85��GE�	�e/m�vG*�$!C0{�CrxDC""��W8�|S�/�O.B���PY� Y�b�rzC��6^LA=����鎠�T����ph���f
�b[����#H��-\��R�Pd��䞋GD��4����,ݚl3H�$2�_cLu�����W��h�ֽQ���+��@d�#�;�i!̾�s��8��zwꍺ ?95��M�#?G�%�NJ��4ӠR���۳R�bS�F�*�&C+��I*ؤP�;�&�&�*-!�/��/hz��b�:�F�ܸ%?����m�&<��@��s6�*C���	���QY�>u��� D_<)�tYXb?�ZA������Qz���}:��ǗI棊D�Y�3��dC.����9��#VI5��������W?���RFRq�P�|-�%	d�B���n����M�0�-�CQGO "�)T�#������dgG����'���R/��_`���>�f���^��g�1m�'�,/xZ�pU��l/��q3��ܲ/Z&�7��f-�*�u�������pg|�ꌅB��H�j���ѣ�[�Mȓ~�Ȧ� ���2f�XӀǩ��As��J ŝ:&?����}�����G�t|XN�5�z��鶸�Z�3�葬���&{�/L]�����2���8�۲6�]+�L�kX6�g'�����qS7��s�Er��g�c@әt8��V��p�-J�`R�z��M}��ӂ�}fކ�J?Z�b���DR5R��vV�V0y�jbY���ծ@����G��)a�:�s�W�i�Q�mn)Wu߂
�
�(+����E`�=9F�m�~�E� �sKs���;kYk���0�"?�c��M�t�`3��H}���w���2ND����4Iq^@�c>���c��
_s]L鋒�o�y�E�����hi�=��A%��/v�����8F���NW��1#�\���^S�Ͱ��+/�VO�'�i���6��g�+�y,��_P�J0�Vvh%5��j��L͔2i�Y�LN��ö���]ຶ{�0h�r6l�h��}�_)�*�^�����U�gt�?.�U�A7W���v.e�C-�Lc��ēT*G�\��(}��r�� lя����q�:�`DA�=}�XAjeV��V���]���p����W4$��jK���q�s+�LW���W�|�5O�?TD�¸�B`����s��$��-������]�'�f
.���>96��j��4�¯�������gf�M��@�r�y_�:&(��}	���C�g��tDz�H�����M"5��	���Ra�s�w�=՜�Mɖ�řr))�5&�R�ZH�0��\S�Y o=��x���H����p>��$�4��H��mtP�zG`��Z�ތ� `>}��&�%/DH�Y�@���q��]{�&�KQ���\���g��2��=�bk0˷��I75q�ϔ^*{�6�c���W���j{��:����t\��V�(v�R�SX�����"�aU,��?�/�����
�le�e�X�r]� ] 5�Y`¼!���Tf�sL�c��M��0���\��X�<%[۞�1<Ϋ'�b��&w��H��w` K;E�T��_�	��ۖ);U_��t��b�����bKL��Jj_qZ)"�>R1���[ceB �v-�a�Йj���u���!�g��]���{]L?��`�$��nzd0טD�B���^��n�Z�8u��ۍ��g��������Qڨυ[�_�Q,a��E�S�I3m�ߠ������(���f"����� ��ƕ,\���Xr�[��!�7 �CM���ך]�j_qǡČ�����[�ߐ�C�=��nա&�F��~|�� �D�p�GX�ײF)ڒ��s����.a���t���O��Y.}�Ⱦ!ߑ����We���0����UY��wuE�g��?��:�Xc]l��'c�/H-��ksQ���������ȳ��_�5���-���136�E�g:pE@��Ӆdb��^,�Z�כ�t)#�%C�OdKز-����;��"�z�zU%�z�*u�V�}!F��t�ҸPb��w����ת�ȩ��-|��%J,�h�(�'VxP �kb��ƅ'W��ۭ�,�I�`_t^2if*ց&�;	�����d�����r6��z@k��gz�(���LoFog=�\~�݈������c�"��^z!B��9N���i�t�a��,�8�H�ȫ}-DՍ���:�:�'�P�+�Q��.�1<@o�"q�� �L�����̲��Q䄾%$;a��)o��eׂX����f^�,�5Z7N6]��2"��;6���� ɥe�	gd���{\N�����-Y�Xu�b�\���E����v$�+@sn>զ�D��k�A�,�w\8{yx�*�Q<`�����E��`��Xj�Wl7��S�Y�sh�E�&T���i/:Ʈ�:�?��
mK&��r�<)ꮣC��_�Bm9UgwTd�u	�Λ�F��e4�y�:�T�Ơ��>�&Tvd��v�*#�:��m��N�GO����Fz�Pm3<�{:�:�KM+t�����9�.����]�����>v���<t�}8$��R�"4z��9=�V$��6�qҊ|�-�����;k`��,KZ�Ȣ��|kD�)d�����Z�x�]�`�ZcL�U��j�[UU��["��K3�{A؝�tg	�����s˩���L�1�8�X���x1c؅�tP1n�8v���N|���H2gz�T��싼�_���X����>l蝍z޲ �� \�f�}{����}�"��-�08��7V8�'�����ʜ@�*��5(G��Y7-x'��B({�u��T��-v:�ѽ����+��IX��a.�TW��ٚ�I��w.�tx��je3*]�F1p��J��)RT���k$�W�6��;X�i��Q�}`����,W3_7f��>����!���a��E2T�/�f��Fy>�o�YG��1��$&����%����1~vb��]�&��>{k{Y���;a�>��VǏ��d�/����2�_�u��n�e�jN2� �֖�2A�]u%!����K;���^�>�F���I["�衳5�����D����	��[���B@��wu±~��yBܨ	��娀�g8#u*�Ϧa�ɟ��4�=�+�
R�Q^[��=��a���14B���G�v5��G��-�B4q۸,��t�@�u'||bD�ԞO�O���ڂY�H�`�L�%mJ������uا(z�Q*K���@�S�Bij��1����m�œ��+�HG6?�UaA��̚+<�׹^�Ќ�S��͎>k�*��ݷ]z��ߴ�Z�}�ķ��=�@l�I�vS��)������.]*�j�Ɨ%Ĵê���y�zC�]p�p~p��0BB^�q@�iy�-ƗD�[z�j48l��[|ì&i;cn���F��;�@fw��^���p���k�0=��cZ݄ �ґ`�a=R5�B�K���(D-s�*���G���+.!�/z�SiF����=�9�%�F�e+����46ӵ���^���*�"�nd��@%E�Š�����"�8R$UY�,�"(e�_�gX�<���gDpf�������;;V�UL�z2����QF��M�Ҫw@�0�o���C�R�i#�r>�k�/HT�l�ޏ��!=�*܋� ���Y������&��u'!��N~&��0&&�D�|��ѡ�0q[gm��:��3��������Gs� [|}~�W�? ��U�����~ZV�E�l�NԋA&/P��{��*�>6�M������𾜥�9kB�	��!;l����5t(���xĽMt���L��]�ŧi�}'��j`�Nꞡ����I)�/E	������y�����Z2�����Ea;��ۡ���	GW\nG~>fؓ�X:gv�����Vۓ�-~�"�|o@ˑez=ԍx��2��D�-�o�J����i��EZ�޳���̸�
�q�P=���T�f�<؆P��14�Fy��5 W}EY�}����]UR�c�U�u�C�^���������q+b5��b���n���ʔ�z*����������r�ОhJ8�3��d�'ة�aY(�m��I>@�uk<�>�ɞ��}���<��&z�p���"j��O�<i����u�Y�;�F]���M4N2�qa�#b:�i�.E�7��tL���Ƕ�v�z=����s�
U��C�U�9�Wڃ�*���c�%U5u��R@`b���^r�nQS`�s��oA��X��U6��5�)���\��[&S��a�H�MʷL:@�r\����u��	>ػW�����,T�52���YFy?�|X�K9{�4=��!޽���;��y8ls�Q��ά�ro����=^CT���Xɹ�]�3�oۓ`" ,��_��Q�(}%�q�Ӗ��;9%v}�2+;��)$lJ�Y�*j���b��_~��%cx�1�?-�M�Wh}:tN4j.�h�2g����k>�X� ��-���>n[0uа���w��?N�{���M6����Bl��sج����ת���q�%�=F�8v�����C��?Pq}+,9Nq1�.8����җa�� �@N����ϩ�wXS|�䇉՞o��oeݙ̻��y)��H�/w�z�
Ґ��l�c������l:�|N�������xQn ���3ɽ�ɠ�i0�&��f&č�����XzKȇ�&���Xz���c^a�Ko���I��Xϕʇ��?�^�B�^�[��`Ü�4�o��0L��+7� ٙG�p�/"^������y6�m�l�	S'ީˡ��&Xj^S�8������)I~�n�ٲ�g��j�?�r�>�뭹6p��&v-CJ��5��4>���B�2��G�}˶�%�,Q�{CD�gN)"�I����(G��#��eTld�fN㼝���@�كo<����7G �x� -f
�Q7�FЀ���ck���)
8ocN�I��yp���O
�(���V �GQG��v�9��F7�xj�N�zs�p�+�V�W�V+�,&-�@��wˏw&��H}C�X@��c�{�b�)	Z�ye�!~{NX�ԅ1(�3vؚۤc�Z))�!+.U�C�rS�2|[��ٮ�������b[�L�M9�8�j�Ǩ��VR��i��[���6�H5��N�y;�w3��縨�Q�;���9c�B���UD��L�+��'�"����]�ʋ���*?X.
�b�����*��m��F�QV���\f���IX�٣$@��7$���p�k�L0�����ղ��׸Σ�0�)�?\/��-��h,�F�`pj�)���l�G�	)����]��i�*����F�K�}9��-!��&�W�|M������}�P44pҫ
S�<��ð���]�۾���9�]E��Y�˕�)&���j��`����3a�+� ��*���&�X������?�00Q�`-�0c{�8�%�33^_���tjL���Z��s������j-�e��g�*c�Ie�[b�A{�ɳM��:=���`\'���?��!К�㯆�g��ǈg�@2����9�#�����Q��N��K�������(+ ��� �͂˩od�����/��0(Ϣf�y�ӷ��r��ZwU\w4`��Ҷ��XP˾��gӧ#ݕ���J��@l%�΀QX��-�/��1M�S��'t"A�T8D�P��b�9�u��ȇ�P0j""�r]���u��,v�$�����|��W�j�ϒК�T�,���2ݧ��/9�Ys�V�7��v�GR3�ܧ�o�BvN�C~78"+=Z�2<ټ[�8hҗ���- ʸ����:uߚz�0�==EI��Y�U[����`yiR(-��ٸZ�.g��^��?��3��F�U�ѹ6[T�y�`f����q�3q0�����Kjcޟ�b����a@������m������s�@$�ӘX1�3�Sh�z�D�����v�Y|��9l"��*�TS��'��ꦟ*��k�D܋���<:٤�=[Y�&��M���yA�s�缍�ˉYP���h=���|I������2:]�ח��E"��O[�~4>�*V�����1tw�?��w9��p�O���?}�SȔ�(�x���##�U���gY��������j۴�WV�{_Ew��ھ�\q8��8�Q�Jp�P��|���3�d�K6'�D�_V�W�S�ӽfŽv�i���ܟԦ���S%��a��'=��F��	���,J����|�5�4�դ}��x��-�6f�[-���7��m�������sq�K��R�T�N���W�a�L�7���E�Ed�S+���@�ʑ@*���'r�,��v+�"d�B�:����i�A��8��F����oQ_�e������K����yq��n������7�<���v�E,���/�4Q6u��̫\%yS�	�rqʁ� |t��Cy�/�IG�~����L� ",rVwȣ�"0J��/�]��Y:�9�+|��N���>���%�z6,���LT�*"��@d��u�L�;�?=J6�GX�P/O�>�`����pfȋ�����Q�0i���9������B��z��c����.�M[ަ���i�<�w�R7%n��� �/9��RX�@:|�po��dWѠ�7b��`rB�}��/��
ΖP�e��V�}������g�GV����~!$�k�"Q.���c��Lڰ���+6����+�/.S��]�T�vB'��V���8��ϡ�0�(��_��x��7H2��r͸#j��mB\y���'<�0��?*��6Ij� dГ�_�t�c����M�g���⟰����3�)�>���E�J��~��9n<w����m.R�����2�#��bz��-z���L4B�7N,������2�]ѩ��=�j)���
��G��c
��h�Ł~k�{���!������p��S��L�o�	�s��Whk�>x@�Vս�����qh���a��&���� ���^��i����-���l3�ꂟ=�M�o��f��܇Р��T^��_�W7��&<��M/�z'�d�Fs^پ��3�i��A�
`��<�c�1�!#?@l�D��XͮVy�DIf�3�?����Z����R���/�N�-|����C�K���XYu�O�Z^�Il���0��t���s�S�����YLm`����p%���}o�գ� ����I��$���5�@��A��,q�H��b��c���zw�u�� G���B7cj��¡�O�'8(-`���p;W�,6��v8u(�U�)��ܩ��Ԡ�}}lgV�oRW�g���"Վ�M��<bG�
�-FSIYF�O����Cf͍�A�J��U��_VPM���bsxզ�����5B�ˢ�t$O�Sό�p�m���#S|;��q�&:B� ����q�}=]��<\����3��:��,��b��ߗ�B������tT�S��gsK�].�5�T�/j��F��˘���q�	�A�����'��=̓�c}����Xߨ����Ob5O��6�VDp�g1����_�y�n��*A����#���ߴ~�7�6ҫ�W�Ր��
 ��Q���~q�' ٪�F�����v�M�a)ٸ�ݸ�q�Do��ml_��If��ߑ%5���C�3u��CS�
��97�������X�
!�ꘌ>��@�[�aZe���K�>���_�E���޻�7.A���@S�j��!�QBX�]�}�s ���s�<
V����y�±�`�9a�$�(-�8���������M ���h�M=(:�����N�c�,ɷ�ޯ���L�A�����R����>=*�U�c� �����P���>X����UY��W�w���a�πY�K��J쥈gCfv��2~F�a��B"��16�������)'Q]�"#6����'�P��l5�=���lQ`/��T����~k��e�I�)y4.<��>����5�*�8Y@P�`�,Qr�S�ʂNL:v��\s�N��1��'��w�n��^4m�EЎ��_���:N�8����(���h[�5Q+�t:M����'9d���X��m�\��KX��/S�\�9.��6tl�v��TM��bkm������C<Q�~8��z�������6�9�ڻ
1�rPRԧ��� ��}_��c���mqu��kP��1�kz�aYgڣ:�v
tA��A�`�n��h,t&Pw���N�ݠ<3���j�,��._�����W5�T �V-�[��㞘���N�]�-5hb�M�s	>���}�@�}��z��>�ޔ�ޓ t����җBcj�{/�,�}B��³N��	����ƽ*�c��\�qj��Q�	������n����w��0�.�~�^��p}��F���J�Kȶ٢p�YD�c?�z*��9���]��Ix�1��ztseuTZJG�ŽC�F���$x�Y�� fbK���i���P{.��,�w�P}
	������E�_��Y�k@�T�Rͬ��sz
����:¬'�xwdvF��e9=2�s���2P����z�����`OA&b�4��KFp�,c��^f ��r婑@K*����i+���o���	-�SͱT3a�Xr1�&7Zr�Ol |��\�&�VdwL(x�w�i��X�&��v����D2�l������>�K������$l'�|��k�eVNmz)1����@~b�WGhJi�@���W�����([b��,#c�� �j���'���g<Q�2ZTM���'8t�l�/:�¶�����XJ9��̪�A;�� �Gd�w�
�/�f,/由�AsnLJ��*��Rr�<nڧ"E�3_�hb����Q�ү�6�R���0�2Z�8i^,������%Te�V�A��~s8�^�Yg�P�0�g �_T�1�tۃ���(�r�!�½�U�U(3��R�xk��-/���%�RQ���v0н����'�?�K:��;�xS�+��<����S	�����&���2�k��<dr�`�%��о���3̟Ojhf���}&1«�"���I�{�$O�<�7Xˑ騣�|��4����D-�a�ɋ�����L {�u��,�Nkq�L*d!�;6Ѥcu�Y�w=��ou�"�H�7id�,b�̘�[=�$��IU}
J׋�P�6u�AmO��;���L�X6����Ȝ}!�#��P�2����#a��ǧs�4!�.Yr���'�"���ͩ�<7�� kl��
�{e�$|�ź=ZAK���n�E��ca"x~�����,�������?d��T�ګ��Nܕ�Ϋ>��4��3�l�S?���	����o�G���1�s3�a���L�T�x���x*D��v��~��!�2y���'}M��v[����}Ht�2�h�;�+I��1�Q�}�4�q-�uX�]��ϕ^j����������U�q8-���X��(q���D�Ȗ2��{\�)Yn� ߩ��ß�$��ʘ�`H� �~���P$�B���m��'z�rL�Op�f���Qq�W%�S�1���yϖe]+���XO)I��ގ�p?>MmZh���/���~���M�6�^�����x{��l�?yn�lF_Y��,�n�d+���e3k�~2&����]]�@F�r��w�kr8�,�9:�L�h��6pR�C�3���ĺ2�����ꩻ
	��夙�ҧ=���d�IZ
��޹.��Y2�{؀�e]�gV����$�p���\4���8��t��Cj�m���%[cS�?��T�##�{�H?�St��%��[}
�f�蟉������@,�A1�	�"^;���x8�}4��@�3���{1
,��0̖�*/�B�g�l����Nt���Հ�!������G[q����w	f8��k�, ��ݔ
1&�C��;����*�{K'��/�a�������g��3��H{���U)����T=�>.D)�Lj�-?U�[��,!�W�<��ɣ6ۣ�2P��&��y��;�x�C�{h�l�f���m�~�M�9�W	w?�d/xI⅐'v,���"�
I�\ꋃs�0���H~*�f��������~�띇P&��:�*��@}4��B���
n�[%pZ�Լ
Q��������E4dTy��P�`}�-�1����e����uo�.�)�9G��r�u>?��]B�[�	�1�n��a��(�s �D"�oH����Q������E��[ 4�e�`d�u���8����ӓ�"s1�7V�=L�b�8�d�Wk�e��s��ܑm�����|���B��#�7"�P�Z������'���ջ�>�K�tL�;�����́d�/$�Vi{U	�s����&{F��cZ	2Ð
�o�-�У]0)Y�t����Bx6	�<�u�Oh����U�X?��5�FXQ3�_%Kp�S
N��7SZR�W��n��&b� 	���~ѷ,�aIp�7�$w+�ʜ�x���eΨ�R��N6�
[M��� 7��mI/�N�
Q��n=��ܝvkZ3�jݠ�`�H���&#�p�C�;Ո�LZҖ��F`+K7^4.���~䠢�t�|4�6�/�i���f�p� �t����+�$4m-�U|�4��]�םťm3�m!&�1�S|+�C�=Ag�죜Q����q�z e��BH{G�e�3�����f�-����t#�����S!�����yY˼u<�w�kn�����8���l�ʺ���V&7�ӟVU������`$m:��O��+��-��${����\uh���`fѣ����F�`�砋���D72l�J�s?��d��C�.�n�`>��h�gnfD�!т��N�L��6�l���1��# 8������������1Pi��6��!�ܱϭ˼m�|�C���
�_0�s_�~t?(ɼL�M�b*L��w [�"������87jA#���?���8'}�a��sg�s�C?����T�lbpdd�;����p��	�����8El{$�_g<�ܾ@��,M���{hNX|#7��Ğ�i��@�}�_+^��ԋUV�<�7>p�_��˹R��΢=a�����=�z�Q�l}0�.v��z�}=��b�[^���"Wm�%���aGd屩�Y�TF��*3�rB�E��*��L�fجs5
���eZj�A���P�a���6����׾��m��?֟�d��� Ⱥh8��r,�����y�J��L���������m��,�Zɰ��
<���":0t;������29�3Y����)�ڢ;�T�0�-Be� l6~7MZ�UB������ң=��h�s��G�Ap��x���c��Xm�%��Ɛ@�ЎXLo��6ǡO�*zg�m��<�f��Ŗ��X ��T ��m�\��^gf_C�`9ю
���q���w� ._|j\'�N�r@,�6��-���>����7��.�U�P�@�H�=��Шa���^���N�A�S�����C��֘Pt<��jB'U ����Ӓ?�E�"djsM�X%� w���)^Ma���<zP�JP]pp�et�_p��H�xlͰk  �f����U��������5ɱ���m�W�t �Y�G��N���'��r��Hx>���������ć�J�����Z3��2h'�E�\����^��@����*��e�Eܪo�A���w?�Ή�C:���<�3;	Wa�O���ݕ���?�dm���R����<�=�,��h�{!UҸ����[;�_���%;���`6{��kAG��LD���[�?��5<T�����8��:؟!�8VRg��MΑ�k�o��;Z�UƢ��i��/�����JP:�v�C��g)�Fl'�-R��~�j�����lz邥�+��VEQ
���!sǴ�9�4� C��kh����:��Tb��E$�P� L��"����gOL��BV��Z@�4������6u��[g=�D��D�D<�1^�Ɋ�M�#AsIJ�EsDN�Ş���f)�ݕJ���Pړd�`Щ�n��]OO�U���*J^��>RGz(�ㆰ}��t�<gW��Ǔ��į���m��5Ig#��q@\rMc�!��\Y����s��=y��2�{��n|�, ���q�Y
���(�4w��u�p���I��QG"���6C����p�J��hL ����xT�� 	��x���J�w�DW�HC�XD��v}"�s�t� ��iMe�{���c�ӓ`�����.�#�zJ�$/yj7�3�Sp+-��B�O�.."���;S2hi�1�\J�bb
�!TV�}u�xt�4�Ki�x�X�ɽ?��&�]�н�#GP��w��U��9��sYuR����)xy���#_VN��+U��H4�a��>�(
��S+�H��k��bj�N[�u�69��Vd�Yb&J�ݭXY	�$�_#�r�QY��eW���s�|�ONĎ�����DBd�
�z�<h����ߺUJl]�:.�x��b~)�g�cO �<xP����٣�V�a��h𑂨j�\ځ��yB�����9ո2�Xf"�`Y�Β�g]۸�:PҲ7nכV(4��֝;��!��PY�7U�Rk���h���ka�`�l��\T�W���:��
/���,�������ݥ�oI�9d�	�dz�R+m����nr��j9�5�S
ъ��M�v���I���6�%N���'ƒ�;}q'��cUxh��yn���HO� Ң&:��� j�?��[˂y��d�N�Y�8Ht_��:�h�nbo����娴��T7�W�&s�\��ȴ	c�ԕ�L� �N ]�� .ꂄDr��ª��{*��i[#Q��������n-{}�K��ز��5%�O\g�,`896Z��㱯�Cѩ&�5^���Z��Y�4ƎH����iV���HD��]�mR��?��ڠ�y���bH���(5�	��P#�NY��b�[܃os�!!F`�㲶��'�o(� ��&�GP��ӕ�4�GL���}6۰T�-;x�|��H�d�j���������A~1b �>��}����u��$��
�5�kLw��qP��}�	���z̼��+?1�,��~���Y����~>�1$7t�9����͉	��?ًPzW����V��8�g9���Yr��`����y2A�y7���Ξ�&}��Oo8(�~w���]D��j�#dAc��|#u�c΂ga��gÁl���+x�qz27��`�HR�
4�~I��HkW��u�6�I/K���HA�3��-@]�)k ��+~�M�EԌzl��/�r?-c��Ci/����g�* �Z���ͺ�Z�iS�!`<����ֶHP�P섒�\vS���"�}�+5��=�`s����h����3$?7u���5S��"�Sf�Zu��OI^&{����/���oc�a��u�R��M�K��L���<N�D�4e�?��6������jR%�22�{v���N�f�G�(�w�FP�s}_n�=S�H8��_�O#��*B��`�O3�ID�ў#��������?J�#&,�iU�Ao��ݜt��%�v�h9n5]�s+2cp�d�hY�dt���>;�+�����&�3��[�wT~v20Ǖ�ELjE��Q[�R�e�����[�h���� .�sMZ�d!]�K��̮��V�6���2)�B�����hDm�=�M�Ej+G�DP�r��9N�7xI1����R�%�~����Ti8���_+�x�X�/y�Q���ވ�Y�B;�-ƒ]�WR�v�]Y=��o��ˊ�{�l���:�z#>��0M�q]nfBS��X*=�u&�>�eStw�u���+=ܕ�� k�a�*~�ktt����W������RЛ�G���m��;�$pR�W�`����Y����/��l��PG����#s3Ԫ�am6T�-ν�W%ev�!C��k�����;��V���T����<Ό����U�K��� O�,%+b��Ҝ����M|�����X�׿櫗�.���k��R�"V#�&��LH(��lӘ�;cx��_K�v�aY��r6t�]#�,�ƯsWt��1"����u=��� �|J>����&�I���˲,����n��_K�A�X�E�-�|��wo��5'4Ut��2B{���\y�[����lp�@�aj�d���:�Aa�H$���B󨙿<ڎ��vk�#pC�[x:IQ@EI<��=L�8����>1��F�ݶT���A���f�*&G�}��' ��2�i��!��X=#�up�tힸ��FL-i`�4[��� ��Ĺ��n�mOAzSY�?�;�W��������7Б�ǀoJL������4E2�����|)��������O�����>��#�	R (չU�K�)����<Ѐ��|���p�DY^l��� ���0�8�������
0�D�����$�|r"g�H�/`?q��"�ey���g.��vs_�7�@�q2K�-˳���;� k���c���5$�"����m���dd�G��g���Z�<��ST�5��C�M��Ф���DEq���*?c�LQ�_�����̾���;f��3]Q�;(�]���D���,%���C�5�-���\�r�1���k%���1f<Q����3h�?�E��@�8C��!�D���1���IQm��3��8EY��;�ޅ�7z5Hf(�5�%����$����\O4�Q���y�#kB�3g*�LVW���ze�GB�S����rL%���Ȓ\!��m�d�Ej2��ea��5[u��9C� ��wu�Ǫ�6���P�^�Snd��vFB'�L�<�2 �;�������)\7���Y�O�t���G�����ބ����^���R��{I����*n�����^���uջõ�:�­��[V�s���?���DTr���j-��i��cXI��=�&
;/�5RQ���0<�C��-+
[i��2
�qW��<�{��`�v~\�+N[~X�ť�+�0�[�G�w^�3���=���GL�Y�n���w"�7�>��F�1�@a�V��ن~�|Z��[�<�g����J
̮�[�=;x@��F����eY���_yхˮQ�"j����O���+V���,�̳`d�|\�,�c��ry�g��=�O;�o%�̌�<���e�Np�d_� �t'_yP�U�H�g�/A0{�A�O�C�Ϟ�`�ӄF���`�Qe��ZS��1T��qJ%m�<��{O9[�@&�����K�.����D�[�V���W����d���Z@F��+�j/[�K:���{�0��m �N�C�f8�T��Ø�r��TK��p՛�e.ݫ �Y������Q�=X\)/@�P�t9DO���ķ�I�ݵ�i=���HA��(�%+�����;,PWe]-����e��� �f�w 	��|��q�4� -E!!��Ŭ�"��f����Ymg��4
P��xN���=������a獺���jB˔���1_�J�g>���$�f�m������@�h@��t�?� �b��Jqzl�w�uC�,Ŧ?��4v�࠾v.?�+�b�xRmiL�B�=
Z�8�mҊ��m�Zh��_!�rF� Y��i�Z�\7�Y�W?���וh�m��(2!�Fm��T����m���Z���S�m������9~��OKp[��I���XG��R-� ��+@�̬u���̀Vcor���m�������ta��:�6}�?S��V��m�sc�W_�r��P�`��y9���}Se�̄Ϩ��W���['���FzDD�K}'�w���嚅�؎x?����tyׇs���nPmGl.$lA���U�?�M��<��p��
yTb5��$J����v�ߦI!�r��3���[���7`9z��Q��[/�u�0���k92q��:�	���P�h{z"��N�g�;ĵ�P��-�YRA�ވ���]h��d��w�Vt9Z�]
�$	ޔa�Z��<8l���>�ô�v�����nm�5=	g9t��\+w6>�`%����9g�k�'��B(YSu?�=���n�C���G�E��h��x�Mn2��e�rL�c�z���0V���l�(��tmi
��� E
M�8���ڲ�.���V�@>���,Ms��hv,R��wvC���!���L���K�t�n�Fk�]���!�����??����t�2p:�g����)�R�c͢�,��Byʋ���$!Hs6#1k���V�R~�[��e��aaN�/{J�Lr��	;�<6[e���s`N��9(�y�}vuaf���l/�%׆�D��麅\;����*w�=9�R�3��Kq���fd�mn) ���+8��{,S�l����YwN�I�S�)�@�R3�0�VY#�yM/>F�z�e���M�Q��~\��@��׎d� /�w�W��Y9mL��0'"��ҩ$���6Ŧ���8���Hx������P�~x�]��8�+��U[��1�6��Un��kj��=8�`���)):~�{*LE�a7�g]��#_[au���מ��ٕ��*�ɯ�[��I6��O��uu&��|����Ĺ֐�i{�/^pm��3��M�W�Ɣ�i�.Gd�sI�L"Y���7���t%V�����Ji�4ȭ�
0��-��߭�DC����V�-%��X�6wey����N�2��fN܊�O�n�(A�<K�ߓ{�r�bG�Z�+(}�d��0���M桌��1���@�� ����¶@7,G�!�i]�0�������8⟔�:�������od�?��{0wg'j�ٜ�_�
U���ԑ��5:&^Ҭ)��  �Õ/���O���T�=/�o�R|'iٺ�>�Jد��u�7�z� �@�g�]D�q�Ψa�2{�`�j�MF�n�m&�M_���n�w��$D�?*�d/,ҧIfO�,2>���.�3!.�>ڒ����$U�
u�p���OT8b�,�P�R��[sZ�1N�j$!_Hr$��*n���[�0`M��k��˜0����7y��wڄ �+ك��#���q"������d��BS�_H<�C O���z)0<6��<'Ή�E��c����R4������i&#���K"�u�Ma���g�5���*t7,�<�ʹ��Z�� �]˦�AtN6(]�Iժ&KҨ�k&��04��fb�} ~�9�qj^JI�8��X[|`i��D1��B��cGjm�n0>cy�0�-A.𬡠����R���2XO�NR�'GD� ۦ#��d8W�2όL���=-_^���ihhH-y����Q\sCg��j�!��m_!���� ��^�_���$�3�h�>�??�t����V�E�C:��J��Ol�q��F���S��bt9*@dȣ,z�Ypg;m�R7�p�R��T���!t��I��Ez��Z$�����t�^('H�K�9��o�d��I����TZ/�H
�$����`�RF;�\ ��55���APiU˔����K�pWc&QA�mV��v=Ǚ#�@-�G�q��&��l�>ʆ�����#�`�bE
�1����F]��,������Ƶ��xW���R\�]e)�	��Ղ�.��2�.��S�n���&���!b2M�m	t>[���ږ :����D�"t ��9P�䐬6qj�~��y怪���
�U
�(�w��@T7��w�^P�f��ⷭ?�����w��c]���[]��pp9B��Dc�A�"2�ʒ��L/�%4���(���U������٣*BD3ׯjjZ�D׍�9ۆZ{��]��ui;�F*p#��9�x���`$��4&1��҇h$>��,~X�y/�"� Q���+L,>��l�Fw��&�4�t~����t	�����.!�kR�A���nto�1��O���?��V>O�l�K�ׅ��܆`���% 6$�ݿ�$2K!��5m@\.��<�0�F�fĶ���͖�14k�b��NG���V�|�ؚ���Q؉ܺ���)np�E}!�Mɟg'�#�i�����b��yK�$,[������7���t��\��馐6{N�5O�ru
�g0��t����D*�=��^a0�a�f�8��� M��I�D����ŭ���]f;�I3��T ~ܟ�3���yp!� o�����Pă�<OSq|Y	}���i�G�K�|�%n�q�i��n�{��/�xFق��Կ6.|����=�?.�
���4�H*s��4i�+B�{JR�#����~^2�M &�]y���Y��nsr�'2>�q~j����y���E��G:�+h�H��pr'���3Z#����MjN(�hی�x�Gꒄ�I�&L�	�L�O��@t�=��Ț3��ؾb�rVG
ɵĀ{��]� Y���u?4�����Ej����~��u�d��1�*+`���7����(c��$N�af���cO��]c�a p9�̃5o���=ڶ4�p\\>��W�5�f�S9���X>�.��n昮��U-1e�0�.�
�Q/���@��2C�(�a�c�?Ȁ�w�d�~9Z�SǒU3e�\4��V��Y ��? w�Uu�9j܊���ɮ�R�fL��o�X�w�s`u~��~BN;����;8D\�0O�c�V�Mň��7X��/��C��`z L�E�^ԂFw 5XQ{d�}�ҽ��P�IYnڀ�)[�2Ԥ�Ǜ*#n���Lć��Ӻ��%2L��eJ�=�����:G��MxG*�0$l7���\�D����¢Q G��Ų(�MB���i������2��-�x��g�@/9������*Y?r�v5�e�m���Y�Z�����������x�d���.)3r����\�Ci[c���Q��M�U궅&��:B��P�'�Dt�O�r���$��l�M�"1��ɾ�����(�$��ؗR�ԛ��5�љ�v�#���͆>��ȻGu&�]�:��!����U�F �ȏG�� µr�>e>9�YiS�O,�8/J�ĕ�J�|=�+��S����;�Q��?"Y�^)H��f��
�;�'K��	�&���N�l���&�wA��Ia~bVU+�qB0��g�+�}��xC���G%@z135�t��Z�BV|�
��2�ֱ":y'��A�C�<,���P�fU2����&�	�B)�8�,ղ�.T�(TtP!E1��Y�jDx�,��f�2��o�s�Б-��}rk�7�Q�A
!�2�C�d���{�Ǆ��FPF�b!�	1�TvEZ����2�t��h�����S!6��QS���� ��L�IÃ�	��r���CIf��u�+YٰyںsP�*�"u,�S�ƴ-����1�Ǿ\h��%��|��p�a݉U��3M[���n�"�jZ^Xl���8\Q(*��o0��������(k�֗O\^19Tt�˺��Da�N���(��g�� �\��8�
%y�Ħ�p��@��5�	nLm�51h@y�����.m�Z�t�3����t%e/:J�s���>���m�u]�Om&׳b�!W�/��g��y�tgd7�;K3��U�]Y�Gi1|}��z��~��W���Q��1���vwB�3;�^�M���Mݳ��H�aĄ%����\�n�۸	�"f�#�=�G@�ZQŵ��im�+t� ܦ�\����9���p<@]E����shPQ@�'�Ut['*�LJ���BYD@e��U}��pi�6[�g/XB�ZZJ����?���ʟ���o)�B����'"��}��EO䧪 ���)AJI�kx��2�+�S���//űxK>TE>���w�g�s٬n��	[I~t���R&��C�"!q_\	��Uѕ��Q���g`�n��k<�p�����3]Iկ����yx�
�~�R۾N���3����6�g�eUJj��ܲ�Z�n|P�!���ζ8*��� �='�g#�}�ۿ!����3�5��L�hmŴᢖ��q9I�)Ub�vR	�[�Ut��[LgM��W�.�6�� �k��Ф�`���f	��8�q�n��d�N6�f뉐&!�﨣�����������@�g�[|LͿ,HrF��Җ�d��g���F�Ġ�i�.��U�F��~�;)Y^ܙ;*p-�u|9�j�cK���`G[�Q�=(��B[2z�`�2!�F���Mԩ�����#;�V}j1�<�-U܋!�E��׉��&��L�"�����o���
)�JyEw���ܜu�7Q"o�r����������9��c{.N<f���={?�J2l�0/�Lj����"V]p�������I�s��P�ܮ���a�|��u�I�5C�Z�!i��-�G����}U��Lk3���᪳6[kY�o?i�u��^��nڡw�	H���#cn	C�b��䆴*�̆�)W��X���������u@�}P�ܸ�-���pu��.Z涀�a(��4Q?�ī����wu?��B�M�Uࢄb�|G�Q�bd�s�B�e�x��R����KO�YF��3��3�:�$#'M��G�*.���U�c�p���TQ�O��������"�D*�^N�,��ܛ�ma���U�E4}'f:?$. ���yה(b#}��-�9WdΑ�g�LJ��ъ�$���kv�W�?<4+�����`B�zFQ�\>�:t�#��[� x�X� �E�i�j6�z��`����,�5C\� ���	�p�޴K�О�EtNV��F��?�)��X���X�:a�T�Sj��IIˤ}!�����Ǣ���G5�8Pf>a13�Y&#;�ت�DN�cw=��jE�-Ѷs�V	j�T.}4����T�v�]�I�x���{���Z�Bc:�߇�c΀�)��[3;3m�e�|���K���c�����wO�/�M�s��!Pz��Q��95�+T��N��,s�c�%N֐��ʐ�}��v⽕;���GIi�Qء<@�vT	�����@/�������^�$z��}��,�PRY�U޵��ߓ��c
eo6��/J���i�lF�
�� �g��0��	1�m��dhaA$+��Gg�9�A����.����9���� ����3h����<�R��P�b�5.��:E��݈Jx�f���kE�T���,�������K�*�0d!�������X��3Z��J5���K	.u9����݄ԑ�~����$D�{4G�eI�B�x����i�=��3L���x*��X�p�������Y�ڪѫ��瘵<`:�Ph��7gt�� pu߅\�Z�#7B�џ"#O���rX�N؋�*gj8$k$pP�t.�.�^�K��vP[%a�UĲ���63G����U��-Y��yo��?m�q{���~�T���iL ���x�+���}�`R�*����3N$�Ws	N��.�9�C���N�+��o�p)]�Wt�~�8��ÌbԼ䤷�dx)C]	��4dJ�5��'aC�XH��`���ݡ�M���"&��q�q:+�(-c����u�vqm��9�Kq�ۉ��!���7������T�>]�����g�i�n�4#��G�~��t����#��?�i�v�m��YX^��u�ۏ��[C�a�c0k�G�ɻ�@��?ǰxG�=X�ou#oB��g��Ö�K�nˉ��
㶠6S��?�����K�5����a��8d�?;d'٠�4fZl�PӍ'�/W&��8BJ��и�*��7��(� �<�Y����� ]R�l��j(� ��.q\��~�t(Z{Xw�l�X��]��p4�@�H�%s���80�rMisOYR��t�"^���;���� �s�&��&���! 1�� I�PI(��կVߴA�{2}�oWJu] �nlĶ(���ӌ
�b�h�O� �vQ����:�9x'�a�
��P^���E�]M	�����Z��G����s�+�WoT\��π2��lS#�ONVY���ɐ����zpE�$�ŷk��B�b�]>�dÓ�p�F�n�Đ6e4;�J&ẓ�%c�خ*�h�� Ŋ�H㲨�\Q��B;N�e �L���s�j{ɅA�1�8���X#�AN#I�����|��F����C\>q	�3�u̮�k�|��]b\` k<����zf#����څ<y�I�3V\}	�LhΰD���g�117M1�j}]z1���qV�I�O|F6�!�N�'�5��2��a�����s��A���莳�5y7�\6�?\�Δtl��eb��6?�	yw
A�'˃��O(5��?.�fn�h%$��;�~���oR��ةB᙭ti���lb3������&����.^װ٤e��K�΍�}���Ez���Z�S�4')�x�o{D�z�'L=H�ɂ5���Ӣb��V]M����KSh̏�R�~��q�JXxYd����`�xO2&R	3�IAEj|L�6���]A7�������;�]
"�8Rc�)��"9y��v�=G��;�������w�<��ɏ�PD���ljx�O8E�ջ��0�!�"G��z�v����B����۩�7J�sa_�4m	��*w>��&����m,`#��?���1�]�'k�	O"JTP;r����}�\�s*��;Xc7��Q"��?����5`3.DL͔k��1�A��cU�4 ъu%�S��$�	R�. ��~�C�
N��'��;���70��@T=Eu;7[�����+'�H�\����������s9�S�C�S��8��Ԑ����q{s0�bIŧ������x��TN�ʶ�<���������7l/��H�.���Qќ �;����jo=���Bf�|�D�}6��G2S]�zKܢ�Bi���g��n` �$���k�RVA_R��B���1�Tx��ojͼ�@� l̔��Ts
��׺<Ҽ��r!	��Q���y�)}�ĭ�6�]rZo����$.�.H@�Z��׍8����m�ʘ����3�g��#Kmn�Éⷙ�ie�E�U�uu�Kހ�M	�R�wC�����A,�Bl�)���Y!�쥸�Q���+�>��I�nt�l���W�	'y����Q��B���7��F�3=o���,@����8�@�p/�L
B�M�x������\.K�l��v����
_];���R�d�,��Ώ4���?�'�P �8�R��pu��P�t{a��"�ެ�m}�� PB��e}��IG
~���2.Bk�7>�A;�Y�	:��?r��x�X �S6z��o
"�cGO��--v�xHMt���R�/p��a&.�`#�)��Ԅ4T���R��B�8- �\�0���Jf�T(<�$m���x�W#����am��<K	���������G  E�OQ�geB��l_�;��O>6eu�p��P��AH�ǅ�|rV�����1v�6�Y�7%\�X9���* 	ʡ�B��^ܶ��8�Y>��R�0=Ь辇�l@o�?���������q-ɪ�>� ���E?Ǳ�jUs��e��xĳ���#�X�B��U`�������slj*��}����3^�),)/��s`(z�v6�]b͍:}�m�d�U*�Be6i&'�k�c�y��֎2�<ߤbD��[64�aH���᡹X�5E��;'�<8��)s����O0�^Y�����]4��E��1M<5�u�o�����ό��S�[�N�RQ�0(r��M���#�p����0�<�~Ȝ����g��[����׼�Z1�����J�J�JvB���%B#�f��/̂.�$%��V��&�o�kt�!�Ы��{���Ⱦ���#w�";�I����=8/f�ۍ�Ť�h�]���)�]����wiBK�nU��0'K�#�>��^���fܞ���X��,ϣ�	drgZLN��{�Zl�qGE��>І�$�a6�>�E/v�0�q	Y� i�QG�_}�jo�ћ�~�[䫾�[��|���B�������_�"��j	�T�����2�l�Y=���v�12�2ˮd��I�����L��2�@Ϭ��!�O1+H�U��s;�ye/.���k�)s��F�dK?{��
#������'��I�۸���O�Kl|�{��&�]�aA�10sR�B��;αlu�Re�ݙ�e��sǖXk5��	ݫ�����ar�Sfu�v����D�ЀQ���ؘ>]2 o�շ�'`EXn�RR/1X,B�l']o��Qf�,,v�Ϭ��]��wi����>��T/�N�.hNg�����h�?'GuT�<��ӰL���'����d��_��#i��h�@�F�i�caEq?x���q�.��V��]����9���ߺ�X�>�����r=r��s��n��ƭ��mR2LzD?&��:z!^��,�W^�~�U�5�R`������ýG�[@BKμ>���c�-��@��̪��[πy��O��`U���$�tL��sҼl�un�Va-Xa�H���������s��Y����;�I5~�_�\��-����W�u�H:р�zv��.;8r�c�h��f�h�������Bz�[ 2�r��E�5{��u�i0E������u��_-�L�Z-> �p���ui�`�rΣ��&�pTz.��%��/`�~X]a�gb��\!���#ց�1#��]w���B?v�!����r�����>2���[
Kؘ�y����K
�qz�;���Q �m����/�2����.��}W��K�O{E�u�I �*_�<ųⴸ:�T�� yJ@��q�&��禅���>LKQv����9=A|̐�������]Nʗ��`q+س��ĵk�_�u+��U�o:Yo�O���L���G�my���>�7	�B���F~�Q�n����%��kVan��vm̀s_Bu̇<����]Ȕ�P`��E�Ӑ���dh+J��Ez�_��u�e� ͦ��9��t��Wȥ�C���.��R|��u���@�ދ�*%f��<f��-���@\MەK-^�G�.p�D�=a�,:/��?�ޯR0�̶K��R>
�ڤy��UC}>P��ÃzC:B	���&ڟ��t\�[�^*��t+��o�XMF4�~�L<���%�׏	��$}���r�K��-�@:��;��"�З��x��������E�Iy-���~c����a�$�����(|W=�ŉ3�A��M^�&d��=ضĞ�XULjm6�:A+Q~Ǝ�)�`��.6%C�K�lY��*�а�C�F^c�|�Qͼ��,TN�EAi���E!$� `�m��aTN��jh�vd��:��D�b�*�r�����n쬍8&�]^� y�V�/$��:���x3�S*�W�Z����h:`x�*�ӆ�����.S&��^�7�r��oI'x~(�|
}����}��k�Q.��������Y�0�q��GKgK}ܩ��lS�l��_�GYMcXl@��>��?1��_Tz���P����R~�,����u:���>Խ��C�N��L/�4+��1Uǀ��Xk�\�e�=h>R�i���gV.д�p)��B��gw���a&��Q�0i�Y����W1p_�����\��^�A�CƇ+����`=v1���8�2Ǥ��J��; ��Ko2�I��Ý�u��I�$�nMR}v�l��� `q^�
��5u��`�TA�!aii0���|[:&ꮶ�S�+,�-.�������"�q�hl�3���V<��{iw��~
��Q�Gg�GeQ*�so,_K�m�cnwsG`y;�57e�?E!z|����;�y���Yhf����R	�%ո`K�L�=� ����t�Z�$	;�����������g���K�1�'��+\]�"��NE�F�)�P�𷷥]O�)s����1H�WǷ�x���z�"^w֔'Dx�r飤��Dߦ��]�L)@K���e�.v|��vN���צ�E���nC�.u�Y�MNR��\.��̨(�'��%d�:%80a����v���a���}�!�i)L�>o����[�]�?6a�kv���v�-q�����d/�0��-q���z���:��iʓ�9����iPć���T	����r�� ���X�3�&��r��vŮ�]+�s"K���~�f=��59�r�������1�;<��B��i�F;��^���l���@u��d����{}�~�o5�GfʎӲ �#B���f'�~�ä��_�y%�ż}=C"P$�����Q_�[�9&�
��f�T�Ƚ<���H���@�Eط#7�kADQ����$���#�ʏT{�E����8�x�Oǣ���4^D
����ڌa� �Z˼v�.PG@ދ8���[B4̌�iR�.O�P��K�an��o,�P�v�:�y��K{�)�A2� 7ƚ�E�͎�f��;��r"s�ɹX~4i��ǥ�)�?">{����P�E>t�����\�����6@�!�g�k���@�g���{P�dY�^Hq�Ҵa�g�0l����֟�3�f�}��F��'� `�"CJp�� ��#KU�D�MiM���J��t�s?ð�`�X.�X	eN����Ny�zI�+�3�2%��=\tq2���1�Ǣ��;�DDM��ѽ7��o��=�	�~�&�m�(�&�UZ��®�4�>�.a�B���^�z%q�$sz��Y�/1` �΁��s�V��c���$�lW_�Ql�Q�i#1pB#���E��A��q�A�D(W�7�>.�ř�F��	�N-�*���2)�ػ���3Tg1\'x�[M��ݑx�O�kl��e~�+X649��6��I.��).��@�)Q�
R���/^���?Umf�_MO��J��e��޷5��Չ_�s���$�ɀ���R���n9e��g�'w�sծ�z8����u�c����%9�Y�6�o(D���cx�#�1�xAR�ύb����d���Rƹ��%�F��%?�e�^n|���qx�pL�>\;Pfo��Ɇ!M�Qm�XS�B>�P�kfOњ��X)S��2a�р!�J�\<}�k��Bi LG�끻�s����р�ѡ�eW`f-`zߋ����H���?��4*bkFg�g�$���!�L��7zާQ��{аq�Fl9լXʸi6�_B � �%�q�!+ ����/sx�l|#�P��?ٹ��;I�ќ�S8?D:R�b��q��ı7o������ҤJZ#m����\N�ۆ�D�ω߸#��,�sa�1��&���4�صd�����j:^��^����P4���Du4�������x鼓��lXL����s��r\Ȧ�>���^��0���u�/}��F����g;���M�3iۼ�]6�i2owWL-|��4'�tɧ�nŌ����q#�.���~*���q!�0�}��֧���*ܗ�A�@���b�
��Y DE��\����{�~X�(L��R$�(�B�����qV�����3q
ak��_nwyw2GO�tzf���e2��Bh�P���eF�SLb<���v����!�ӱO.�Y����TgEjzeww�'��D���0��xof\�ȱ�C�L��1�}|��,v6^a
�Y2��r���hf�1.���y�����r�����٪��s��1�½qa�bk�+���l]A9m�R��>�$����j���(�Lz�p9/�E�r���ռ�J�@T>5oMp���б6��;�
�[.^�]���W�]��I�֣�r��ȏ1ibe��ν|5<7t�ٙ|�- �C��g4��$ù=�9ԃ�g��&݂%9W�S�[�;2t��l;���lI�������Ag�|��	l�szz�,Ǽ�r�����o���N�O5��i���g��"��x�R�&�T)�sM
��Ӌca<��>ee%��W�YZ���u�*�m��fH�y�#����ӳ- Ą'���%^��Y2G�wp.�[�ą����R� <�j��M�ɤ��F� �d��.,�n�{���[*R�P��|���)M	��[�6	�햠ih#vp�=Qx(_�q�߬��.���%1c�-m4P� <j)�a�'������j��� ̉K�Q�_�	�]Fsv]�C�s�h%i%�|XΞ������!��T�*W{��R.���NT�J��]�Q��� 57Ű�i�s]�={0V��ɐ�2���!��X�n���Y�P����G) k���~��m��܂�r)�ۋ\
fC� �%h������D��K�F.���;�QL��Y�Z���$��Ko"*K����g�x��e�6|J��gJ�������s�?s�G�O� �CFEi���_>l�-mk���,��߭�뒱�m��s0��]Knخ��+T]���x�O��]l�*���1�B�+_ښӺG"ߪK�0v��rB)�]~�Q��.ϓǣm��ƅp�\7�N�?I�>ه����Y�[���n�%H����
B߽��cm��)�=����Ru/F�&�z�Z� ݉[t6��R�-5W,�9�E1c
^�S��3tb��K��or4*�	�d@M�(2��[��L���#��>��μ�d���@��@��φ�k��ͥ�� �b�	��纙~���;�����Uaz�3�W{͈z�c�;Wg��T́&sdA_�kh���׍C����(��`�'>A�7��ʩ�r�2���%kT}��W��9{�/�@K�����/��.�q����E��6��y���R�?�����{��]#��*���IwF�k�����7��E�-����q�`tQ�`?�'92nV�>�ݮ���t4���fp�ښU��;<��P�D��ϑ}����	��6n��ݦ���Yq��>�,���������=W��Ju�E�s(�4��\�]B��TC*�HD�6�SS0�����9�����Qtl%���S������@j�뿟���-@c�9���3��#���Nfbr���SZ�1-�wU��9nl�r�wE�>��h��d�z��X8�f7N9��]��ɠr,S"vU�^@w�f���Н�}.iQ�ݭ$R]�֧�*��M�!r��d��i��32S~)&�o��U���ac�5e>�V��nW!��?�J��g)R(�{�t��ڧ1���=i�l��J%ذ!��,s0����/"��jE���^j��R���YH@��\��r�^�ċ�[�r�G�*i4v���\O��F 6��xڔ��D(�}�6����0��b��89� v?l"��<5}�Z������h��f<P�O�m�R}iu�G������+y��i����S��6p>j�%&����f�@�n����
���}�J4�cZ�<UN@v�cx?�Duo@w�׽]^O��������c������y��­P1����!fvkN�P�9�r���B\$��̀�� 0��|���3o5i�*�{R�IF�o�"��ٱ�^P�����~��q�9����%Bc!��}m)J�Z�6�|�7$��RG���C�m�صC�F������Y=){�4��.��7�g�J��AT�B�B��7V�ǟ�d.�ӀΤ[�����7+5$hy��Bͯz�^(��U� D�m[E��:$��{��CҾ��F�kRX���YVS��%��h�ÎH{'{84~��F����ϓm�c��:�g<�1.�p��L�J2��ǯ���)�����W�5[@��e����;>����|c�Hd9p�pyW��J������nO�~(m��\�{ń�?p�&�I ����*�G�'m�/���M��zq���\r��%"��	��֏�26kr�4�8J،Hbj�aʛ��qn����?gLHfߟ�V��Ju�h,qJsy�(����,��2X��H95�%y��0fNh�t�UP��ޮ�g4	��q_�\`�ށA&B���T��sR0Ǜ}�i�(=PtH�Hk�]'��N�,z�c�#v�d�x@p��������9-�B���b�^��lB��V��U`	V�,�Vpl�_��+�W'�l���ӷ|�D��Bw�8�?+����g,��z�J�� �s0\c��
����^�ǘB���;��ni��3S������y��ݚ.���:,o��rj��7df��0:uZ�)���^���P�DS]����T�0�w� ��Opɰ�9�Yˊ��zAE���c�]�Ԧ�iKz��y��8�r�%�!T�����3��m�z�D��������P3�������M��T�����b��~��"7�ނ��<��z-�-��<<!��Ǿ�y(5h
��%{ns�́��\&�Z�Rm�]I�f�q�L�S�е^	���������1O;}��y!�s�.zn�C-#>�����S���*2��>�yV,�\ /��Z�@st�n¼ ��'�m�Z�d�IH�b��-�P���!�G8�k���A�������%��%5�&�o��<�g���$}p�~m:��)2�_�B���G	aly�*����.�P��Ь���P����¶9(�T�M����A���K�G-(�E\��(uGq�O3�1)�� �D��)��,�]����R�-)��;�PFW��HI��-'(�cr��@f��AV�<!�8¡���$PP���z:��Y�ad�2]ü�^\�C��ݺ��܍�^D,fMɷ�(	\l�5���ر	Zc�=�qV`��eް�C�%�ńW�T������I/iP5�1ɋ�%�t 
^��6��]���>�E~�k)V��@$}��aB|���Cr�ڈ7��3]����T��nUY���Fx�����������.�P|���{S���`}  ��/�nE��.�"!��/(2����"�.�1��jp:���rf|�
<弔|��U>_ ����ǲ/�($��'?��-x��WY&=o%yS�N�5A�62�]R���9x�56��;M	��c���A�S��(
5�RZ��j�aK ��)W��'?�^Or�7QN���y�"�$2z��ts�2J�r�H�G��;��PB2�p88���<��`�W�a����5�j�A�x�%���0�Fw�u:�8��?:]a�}V�Q�Z���r�`��Zev5���K��^{\�>�P�7�@[}������;�x�c�;�w�nT�D(���.z�`�S�amb���%6�Y�c�_�%���S%�����5a��"J7x�(��%�����C�~��np%���_�/�*+&&�vO!��/��]=UU��������Jౙ��h�L
\����wwiWL�a�9u
+5�0�R� t��1�RhA�w����f�U�8��}�jBA��ߘA�Pq�FH7)y9��Ƴ"#�qp8�N(����:|� =�Fs�g5�c"�1����z� +�@�E�ҾŖ��<���� �ម:�ñ���
� _;khr���n�*a�o8k�B��˜W����xV n�h�c���,mr�E)�8���w��B����x�j�(��Z\�z���_d�P��v�9���M汶c��F�-�&������q/7rQ
���i��_�]$!?����f��,�]���-�|&pa��H (���Ԁ�f��ϖ�P��N@&:^��<*7�.�})�*�����OKg�Js5�*�uP��h��ղ	�Up`�kgXd��	���ͯ)���N���=�0��f� !��8~ID+Eӭ]�U�A���\&WU�̖�;�0���Ȥ��#�b�s0��I��æ�u�����hz$�s�N[oTh�{?P������Tqp�ʥ\��9���q׸�2��#=�'�*I
8�:{#�%�����]�0$��}L�$UBƝ	*��� ������[N]f������3kM+�q����1M��, mI�ynPҁs���X��ĉ8��n�����V1,X�]%�S��>��4俥�h/#����M��y9�'؛{�W%�A��q�����H"h��0�?�R."A���I��sT�4�R�-�Sy� �`R���}�A�·��nEt� �r'}#����Yo[�ԝ���{U�"�]�3�mծ���^j�f��xM�h�Qh�r%S�m��D�X�^�#���g�1~sh�)}�-�"Aj�*�3�J}� #�U��X���w�R��cax��K1dj3��V��`��ғ1u�"���u����`�b�<C��[\>SBF\�6ޙ</�ZV�G��VQ�݊�ʜ��g��y� NŔ��y3�h�f�������9ŗ�_��������:�)�
>ɕ�捧�PR���P�cK=	���Q�ckT�a�n\0����Jm����w'����Z||���Å��������o�jz5F������Íyś���5B�K%�#ٽ4=��������7�Q�~��a�qx�����Jï����A_��ə�q\�˶��+�|I��2��/
?�o[5k�F��������)��f!��>��j&�������C�/�a]��Ei��W�z���s�7:/hU�
&��Q�B������(N#�P}]\���I�)�yw�C�+7`�� �������Uv-Yt>���֤F������R��h��1�ͼ�K%fN�pNum%����'�Q~+�?�Fn:���n�>������fW�3|��3H�L�x
@�]8���j��:w��)v?`��f�̋�����@���m��o<���V&0�O�L)m�!Ԯ�� �	�H�	Y�v�8/e��vb��;��7?c(�"a{@� ɰ˽�oњ�vj<h�f��`�OM���J�a�����݁��9�M�P_,�Ԓ��VS���2�\�b����С̼0N�[Rx�Z*4v���lIMi��,���W�N����T�����=�d蝭�s�s���pث�ܠ6�}��,��.�������<7�N��W6p�_�9�֥��(T�V'�A���c�TZNf�frO��_�FJ�HW& �,�׿������L�R�MY?f�=��9VYvgW��$ݱ*.=*'�V,ҿ���L��Մ�/�<�+��,!X�u���=��=�`�Qn" ��>s:	w`�����#�{�X�!pT�!%Q���|9���Vy�x��4�=>��]�0���m̢�'�&��o_�6�ouʦ�u�@eN��+���IC#�,��
��J������;V���B��<d��~�5M0��:���Y�ݏ�_�'�Ǹ�N��șx�~�U��~3��:�_d�n����Z}����=�rv�~�wE7b�>�3ۘ,�����~9S�@���Q�ˡ��84�S�`�e�߄	f"́�U�W�Y I��@¯�?��+��V4��S3����L����u�д\S2��]2��r%��aOY�>{9���߽�&�(����v�}����zoo�y�P��:Q�ca
��0�˳H��Ν(Awk6J������N�e������L�S��a��3��"7'�!��7�g[�V��R\�f�y�dw���g簸;�Gs�Yҋ��Ɲq�4���  <#��C��P�܋B��	G�$�n+����7���1-檚�,����M�٢u@���k����D�b��p���d0��瓻U6�<>p�eH����C�Y�������g��hf��F���,6�2jJZ���R����`��h�1���xY��áR	QJ�|�.�r���WqF���y���k�^TmRI�����;p�b���.?tO,H�|[�8D���o4m�F0�u�_�B,�s/� ~���	iY�l[C1�]~h���<�G�s��_Q^��w�k���T*@�c���� �'�|^"?����-��"ꚣ�ᮉ :��%?6K�ݸ2�V�c��6;3'pv�����j ��5�����l�%#�\�Zۂ������k�v���(�������Y;���n��R���{��M���XE�M�w;@�:&��]t=���Pc�>F3Ӫn�)�{�X� �g�St�t΃�7�_g�J��VJ�
k���U�y{�	�1�-+�oc�P:&��4a¿��#�^�Z�3���O㥏��s�ɇs�%��|��}�  �����3x����(��ޘ��I����wQ�DVƹ�ƽ'��,��ڄ��=CQ�m��ֹL*āN١��Vȷ.�J�Jv<&�O�mLQלw�f5|�J�Z�>�ET�\��!�GZ�qlw���T8U�5�v_��+_�C��U��Q�wt	$����W�Ġ/�
�ټ�y���%��'A��ȇ47��t^�px8 C����VXeQ����2�fr�F!gJo�Tgt>�lؾ@�k��a�tӁ|�d�l���M���oу�Ҭ��Emײ�}��Tۨ��4T���U4/��
orB�@��d��h����/.A#;D��J�rz��M�!��x���="f�Z�Ӑ����u�Idk�|����������	��C��\J������Ik�V�X���ѣ�mes�_��i��!W����(1?�L~�v��1�9����ەE[�y����uF�5ƴQ��	s��͆���$T|5:e%+`�0�hYh��U�o�=��n�����������1�%��	�\��6'�Oߚ� �:�%hl>�U�qJ{a���#	\�a�I%��ײ`���׼|D	>����(<υ���9���#�����^�����c�X�&d��Ȥ��c�:��VO�i�h�Ӫ���g{�p5?�v$�B�i�g��i�?K� �Ó���|���˛��L]��0�}��A�g	�;��QU������Ri�$��l�xVj��9��a;u���gߩق��B �8u&{fI�����b�a�`�(\D�v���yv�����KT��G=63h�.�D��������I�6֥�N��H#��~z�a�F�����A�T��]n��\O���w�ZF�����E��=�mfQg���ʁX�V�\d�B�^��1�f&�i���_i��wo��xҡq�dٿ�!�f���<�MexCvW6\k:�ҵ�5��.2�����[#dV��}����I>�#ߒ �v�:��
��~��|-;�B2�l�u�Dcf&�q>*����t��s��|O%o���(��T�)M��ED�$?��P����0BK?�Fl8�qj2�d�f�-���Q�ǆ���\l��Lgm����_�C�H/��+�]n��fr5�3���o>'!�mf4o���BG}'jxױ�}3NۻiM,�:\�����`�/^�����
j�ED'H=s>�f��(J�Mb�ve�8[{���s2�w�ƌ\K��g,�e�YQ1wT�^>p��KZkC��7�`-MM'������ʗ��!�e��H�w
3�Y���ܺ.��o�����\�p�"�.iz�L�e�>9{_���VJ�F��� �#K�~6Moҥu��h"���"��������9���o�ɫǅX��(ͮ��Z��"��(.f<l̑�l$�DSS��7q���R�eG� ��NmM��E�A6��h��/�J$l٩� ]t P��l���3�&���ˣT�ι�m�Zl�-9 s hm�US}��Kjڦ�����̉|�SE)p:�TsU��d;v��7��]b����bԠ��4��/H>/-4H[�˄.{�u�����tz'VK[��as�z��)
N�x��|(����=�i��Sd��n��7��ɷ%�J�:s��&G����TWrg�(�8��[�����ku�?F)�ۓ1@�s2�G�&�U �����cS"P�y:��\�OH&��{zr&O�N�Np�q�}Ij��@'��CM0�b2�c<.�����h�]���;R�1?� h�dIIڔ��z��5dmLsp��L���7poeȪ����ߙ�f��'��0���4�����y�T,�G��:��N�3HH��X>۾��Nz}b��'ex���+�eաE@�&��ڷEA����S�D>�
�'�n�Ģ9�~e�Ƥ�>m���7|��/xR��r�U���e�Ś9o�=��g
�g(<4�+�����~�������]��G�hw��X�r�XY�Fols8_Ϳ-��L,Ӕ���'̲����&ՙK���}�h첶��R44��:���^ކO��Ze_��y�H�I�vv��~lH�Ύؕ_��d����i���|��ʵL!b���F^�)/v#IwZd�4v��&��Q�}qs:�� ��Ǉ �_�Qg��o�rN�z@
�I�f��ǰ��U^���)'�%z����ج��p�7�h�X�g��n-h?�V&��O��g$��M7\ �\�x�ʗڿ�BT��@J����ȓam�7 x��뫒��ϽC��K�*��^4o�/'ۺt"�r���(+�8R�c�!� ��myS�0��NM�qE���x�S+ĄF��}���w�Ҭ>G�]
Y^'}�
���q��kWJ�K)6���
�#�������m���ܤTW��P�nB(h�O�N�Wi=�d.�Ϸ7�WEq�nl&��ǲrV(4%"p�a�@|Ĉaэ�̗�<��.-�b�7a�T��N�ȭ"����(�������0�Ź��:T�H�C���MW]~+O�cW$֤�9�W�	��5�X�rʘ(Y���$�>�S��xdA$*���[�7�,�[!�|���1�P���댄�u��Q1[��9zS	�gn`כrR+��}��C��4�!1WYX
���p�ˈ;�DX���K@O�~�Sj�<�r�{]E'�� �P˝��v��_Cs�њ�J��޳i�\�Su��<�"���Z}��T�\r��hT@�d��9eq�k`�٩Y%����D1��.��¹&��R���������`8�в'U�8\��Y��e�����5u� SW�t�5L�xzO�͆TҢ�x�,��ӻ�?���lG";�*L�M�(`u����c��1_�;��-%���%�9np0�-�&� /G{��F5�Q��U.j�يb��U���!s=�T'�J�^�	�*sX��#1�G:�Y�����<zC�CWS�m�k"�|F�Q�'�?�[���@�d#��(��I��*�H�'�5�zX�/3h��,�L�E@��\j	�Щ��3��G8��ĩX|4Q�d 5K,Y�-׊^n\Y��܋�o�(�pM�������O��45+�����!#S�~% c%@��9�<��S`C9!8;\G�J�2���GL�8lZ�ʮQz�����6v�u�x�b��q��M_)��Bȩ8�yH 1�w#Rѝ<��]�U�8Jp�ﯚ�@�&�I	���@�8�������6����nD)���/����q(��K�L��aD)�w�-��_�Lg�v��p\�V�B�eE��������	O��Yw�ͮ=�ރǙ��y�<�0q��B���U����nXz�_����E��gJ��!�f�;�����@T8;�63Q���oae<���/�p_呒x��n�`X����L�V�Y��Y�v�'ұ ���̹��� �u��Uܢ߱B���G���g��)xl���ht��v}]���tDQ���Jv��[0s
�u��pg"�=�l��	�z�J�h�EstCU��#�"�%�WP�$6*.�@]�Ylt�&�H��?����ֻ����S��t^rۺ' ޸.���m0��u[�v�w���G	���o��$���=�'�k ��>&�j��P~���bE�5!�O��@Y2�}���@�f<�T9��s��h�<�-�ν�-����
����*(A���)�i|&�����T���w���M�D���������6�aB{bb����V���;낳n�oK�y�l�Hh�����(��ҙ�uP�đ)])�lH��%�i:S�L�IuI�9C�:��'��-Yn�i�3�'U���|~�G��<���͜LsY����C�F'�Β% Fy�܉�vA�`")?5[����r���h3`!�J��.���8�}���M����~;�GL�W�"��'*ʐEɰ��>�17�X�v��YO�œy|�GL�+�|�K�pEf�:�t7�����\ʮ]�DK\%v�UG.�G��(����WV�7x�*�����{z�o��KG�k|ZGMd��M��f���)�m�%�� �FF�e)���[��(���E���-�Zr���֡é626v�L�ᩡ��dj>@72j�O� ^�<���؟�
��}����=uQ�4���,a�&߁�2����,ؽM!zFD�9�&�	9� 0?�뮂śB��w��ʻ�cL���U��zR��[��X�/��b3��Y��
�0w�r[�QP)���E#�fvrt�S�4���n!K%�C"�F�x�>&)��ZS�YXP��{Y �ʴ��î�b����"�J=�bܟ���L�s�jt�Z�[n�"d������+q~F�����_����+)�
�* �@	l�x����^A��-� p�3�K�ef���%g;�g��|��a�v�i�s9b�Pv��^R�X�o�Y !j�r�n�E��BIV�����G�%ʤd�Ә�H�㢝N�S�t8.��1Lي߸6�W��HG�G���s;F����t��#�W�{(p�2q�(HL1Q��-���[�ռN�ܴ���NRm.�?$���@R��K���y���Vg���t�\�l��~D�H7��(���K����YA�N0�Ag6��M�fߌ�d�͋�V������ҪR�Я������aЖ�3U]�vB8fԲ���_����@)�\l)��<��ۣo��1�r�� 6��O������������$�,Sxh%�T3]��3r��Q=��P�!�z���aF�ն��)���oAY)��$���G&JS?����,$
��_ \�w`(7@ N������L[4�(�4�}ZUk��j�f]߸�?�f��d�w����L{7��;iD��e�����q�m���,�R	R�B<�:XK�������Ң@W�o���\���K{�"�����ev��C��٬�n}: xGś�$���Ni�J���؃K!��?�r5�OCJz�J�����G�wW���{�l����۫$��R�fk�������#�?;�����e�(�Ԕ����g�X�{�G��瓋��͑��z�m��F��(��.{��w,�ⓜ�y[g���x �ݶ�"�|���0���\�X.�Y~�鳧<(�N�������h{a���!A�Mq�Û��t��+ܼ=��Of%<ג���f�Y�\�F�k�;�� ��K@�5P������
`�_���~�>3�� ���M�&�x�Z�M�bG�9�B�HT�x�!fD��H_���B:��B�^{�O� NW�Ph���c��Ǿ¬T����F=�¿��j����&����}�3��΢Ϗ�J8�ȧi ZB��20���Z������������Q�.��q�f��v��o2��5���k-�2<Y~I�:����e-{k`2��%8�N&�z�u���G��9r�Xx�<�8� 7�Nh:+b�@@�B�k�(��F�o�9�Y��R�
�,J.~��6��\/C��m�<�6,���1Ų���0vVܺ�(�T��z��uL�I	&��}TׁR �����4�ى�^���uyj���ͺc��D?���o+l�D��G靈ؽ[���z�Eg���/d�{��tk�#�j�z����V]xj'iK�����*�O6;#,6�;k���9��R��@�k�-mqB�r����r�@?.H��4��$-$}�~��tG�[ww�T��$���O�U#�b������pO?�K C'��I�`�@U%ܨ*�N�/.8�\e���"g����䝨�K��K|���x��+�6$�����^O?P�����q���?3
X�Ӂpi3�x�1g̏b��ټ�6]�9KуU�;�,ǲ4�-ڨ���eg�LA�h!�N�)�����O�OO|��$fb51q����t��-v��^�)�g�Z��U�R6��׆ċ;��	�Y��>�{��ZpО�¤cѳ�j�NgP�JN,�I��R�Z�>#ݴ�_}��a�LS�v��OS�>-8��x t�l?�g`>�HeUd`��ޓv��^J�r��C�NITyI$�
�c��Qx�曲�J�?�Oh��b	���rw�p�M]��D�"Z�!�b�I���Zn��Y��a�_?��Z�%�9�,��&a��:��{�5��U��"l�puW���3������l�.d�����
ZWxY�S��S�<a��"�͉n�0
��*�c�ѵ�1lM�z_'�� ����R��^y��juA��I�_h �{�l49�e�J*\h;�����܇K���	n�����}02˪��o�~�q����9�ɅB�][�Fl}6o�Sl���mu�J���ߣV�W��W%�ՙc`�!�T(��e彘��vtJ��ru�ɚYJ ���ܽ�2sT�R����,���c�0���D��C�	@�Z-�^�u�L��wڋ�G�bqZ�X	R,���J��N��謝����\�U��Y��Qg^:Q^e��$Ҥ�R槮[��la�� �~y1Ƥ SR��Y�NA�҄@+�0��E8��?͞���t�(�63�:6�g��~�+��f�2�"4�<�<�x����0��N�R1�N���I��|*����,�{�#"p����g��S�~K��#7�[��m��Z�f>�K��4H	�v�^_��T���R�v�xo(��l���K��b/N���@�N�^�/[(=��-���BD�S�x�� ���I���Z��l���oA���ڀU��際�n��'mv^�K�2��&邷8��h�sOJ_��'\�os�b��hC�,�1��Q�帋��� C4�p5+�7údDDI+ma0$Wi3�3�������hM��/�o�iaU���i�'X�D��ì�nyĚpu�=��yc&�KG��K�d���������.��յvX�޾������,�3�<��򹘜�W
�ȴ����=��7�~�����c����H�/OP�W�/ڌ�#���<�Ѓ%��t������ЉX�S|�.t���q؇ppX�9-���J�`�h� ���*>Փ��q;�z�ܾ[�~����5�R��B��ܴ���W*����;	R��fl���^z�{����&�
��!��/]�a��TNڰ?=l�Ý:�:���,1l�u�i%��i$4F/?��xF��,�,�~dH(���3a�e��S�n���U"�����-�Or�Mtŀ��(�(��v�,E��{f���6]�1������dA��iW�2�9��6Y�}�H'.?'\��%G�+D��}�4桻߯��VW )���Z� $��h?�a�<ҀԴ(൴'�pp�Z���i�2�$�Ŭ����b� e�3�x�sօ�O�}����n��NZ�u/�����\Ox3��7	�ϐ.x>)��}��	��������pi%���)+f$ߩ-�	�vu޼i5�,���2���w_��GѲ�ʼn&��xԙ�:B����������P�`��8qg��ׯ�_�)p�M��E�:�����h�p�n>y���!*(.�Tq[%�Mb�;2L�-Æ�s��j����<0�B]m�,	֦���D�T�=�Bclg<����3{1�����V���eY�2\�p��n{�ݞl���d�d������y��d�c��h��$�����_���i��MTfKs��{����ElN�q��\������o7}��� p�Y(��5l���.�(�Fش�{Jf�$���c���
%w@��L˞�I��-4��ZpkI��]��4a�3�4�*�ăG�~�N�Nu���}�﹕n�����7N�>�0s�>䢒�V;BD/􀇟��򢏼3X2���g	��8�N�C��ٌ�j�M�X��c��Z0[�S[�Ʌ�K�(����9�����Ζ!e���4�h,���c4����i�� �a
D�c��M�>9j�:R���u�M�m���K4�r�_z�K2B���P�Z:G�z�`���D^��1�.�%��h�#����tjM[���6��C���'Ĵ�I�A���|���B�ܵ��d8G���F�������O\�Q�ϋ�c�&W6���6h^2�UH_�1Vsb�=[��)<
ؓ2������Ρ�<$�l<8aV{�\���7�8!���ڻ�3�а�s*��Ȃ�E#� �����ko�1�8��TU?���K)�T;~���4;ba�u�ؗ|^������W���%;��_p�r'%��ڝ�M6�1������p��
q��c�S��_~����z��j�쑬ha7):���Ρ'8k�j�i��l������m�)�"�%�`=s[���O�� �������Uc�x��m��`RXԆ��e�����-������!��Q����O>k��0�����W�rj�Y�轢���ϙ�N�V�+~ݶ��l��AC�;�v�1Z�}f&G}��bT
>��}?���H�Y'�����~�5�W�>�K�f���˻*��YN\P]/���:#wl͋'���de{�GEG�,�(j'�2�m���a�:J>����Ý�*��-����`����'I��Z���J1��m� �5'�����Vh�xZ��i5'�&G�[bݪ��jI��g.*⡥S�,�vO�Sޠ�+ݣ��t��"�vpl�i�ހX�mn��9�N�����E>R�׵�_�-Zncp�b���-tz��f��
�.��xz�1!�?��T�~g=�C5䛔��t�΀}��)a!�X��"����-�?�sV�:1S�J�Z�B���&����8z:6Qܤ�܂���E��=�
q�?��|��S4JX���]��� �d�%
Е4C�C����i�Zx���By=ׂS����Y/?�(��r�wj�S���`ѝ����vR�׊Vc�'[�+���]h)D|R��(B���P�ECi��Z�;�}_�����a���f�N�"�Ɲc��;Š���BU[op++�:����/�b�#�g>x�gH		�b�����F"3��J�d@���d�E%�N|�ۻ�e7_2�vy�4���5�
&�BӲMk�M�\�SVG�����Ֆ���r3~�b�����E�S	�|�:���7�����s}��+�i��u��-:��6�ڛ�?�"b'�V��*���
���C.�Z׉6s��8�5���uz
"^W��G�fطoZ��,b����6<�̋$?��8q��[�v�p<
q����>�0��*��G|fwDO�0U��3ۉl����΄Xc�5�ʰ<y��GQbtw�~� M2�<	%���"�_���#o*q��U��Ώ�ྼ�%�=X���ʭ��X�țv��oΖ�����B���m������)��\N���(�����t�`C|G����Q�+�Pؒ���пOX�c.��`�����1T2az"}���V��Fƞ�'x�n�)Q�Ɛ*��B��+����@W#{�������K�������D�7��^���P[*p�ɭO��!IP��?|z�-�Fe�U����\��%�^�m�����R����"]�!c���֏�6eiT�/.x����>5)���}�7�%�fizZJ{p4g���[+۪.q�:O2���6��/�]�X�i`"]�w�H�{R�Uo#��p���Ǚ
�uc,��42�vVa��u���)=_=#��;�!����v��E)p���f��]�?.#U���h@��H}{�����Da�c?�aX�vς�a�[����%x�|x��L�+�2]���	�Z�ʖ�
U������es��Rr��c�(��eݣ�7�uLoH/%���i�ˀ�R`���5!��ЛI5������Gd����ŷ2*=R�!?G�\�����7z�*��b��,�MGU��i�����<�|�5�5�x��Uy���N����,�OJ����P5I&���з^SS��/
܍�q�_�IM��훤wa�Ao�,���vB�jN���F����0�o^�U�7X���EhP�QX�qLR^�����j`��o�<����*3A4�/��\���߇B皒��4�h��}�Za�زkÇ�;DA��#��T58K��
�| �B�+^\8�Nq��g��Ũg��'����&&v)-�'������*6�jP���HD�E����nZ�b�VM�^xn���\d�7iGO>��!�ܾ�����c�s�͑�׮��R�!�L���)�Ǚ�c|�g�zS��(�}�������&�3&}�x�J�uh1D����=U��΁��=
���VM�:�iJ}S���5�4,�k���^��s��������
@�Z����M�	�l�C�lö�!��d�W�p�낃��M4�=�mT�t)�,6�v�r�`�X�ap[%'bwR���l�:e@�dX<��tEܯ�.����`�G�5�ý��;�e�	}�|��_��
�f;��k�Ď�$c�<�W�\�ɢH��~��Q^�nc���u�Ҁ=�j�E�L���%B1Td c��G�HM�/Ψbsf���K@~c�y��:d��BkX�'
X�n��i��]�2/�M��4�R{�3���fX�ȭ C���"9qǘ)Rb���� ]n���t���9��U��)���x��D!�76;>��v,�?a�����V�(r���E����ps�v���yZx0�Adc||�^�� �3ǹ�p��N�s��i�Ak��/3Жǵ��)������1K�&x�uS�EFeP>N���?�1���3��io)�iy��X	l�X�m��{�ѐ����)��F9tH���z�%r�����O�&�Z$/I�RsZ/�#�fI�ͅa�񛒵QEL%�xF�Fc�:'�F�W��_<F���D�t�!hXL�e���8���w�A���� �(mw�eqX���J�a�t��J[�d��b&UI7����ɿ�Rw��MJ�W�<	�^��D%,~�b���؏��üA �a�U���E���=#�1�]�,O��I��=T�6�h)/�$��$���Ĝ��K��g���ʍs�-� + ������X�T�G����N
�c~ Sqyx�8��7�i��8!��R9���z \�Y�^�1N��f�:C��D�KU��^i���U։����0��L��tԳ��-N�i�i�wCn�ޫ�Ve ���^`��� �Q�C���/��a��[�Z���6zmZ��?o~�{5��{�L�	���r'j/�ec��C�}����8��"����Ca�;-�b=��ڻ�g#�ω���Q>�6��� S�� W��T��<�ː�PY�����2����!�9��GǠ�w�����C��׎�~�~(j���)���,�%v6�G+���n�q��C�lˏb�ן!Y��Pƍ㜄T��&�'Vd;�TT��QOBU����!�����|�y���]:|����eݾ鶐ȠD����j�.�W俭���e���=l3���J���#yI��3t�����l��(����������G(�;g�!�t��'�qY\�͎�M]��X#?w<�1���4j����Ġ��FE�,�M�$ҥ�o&�`�κ؃��%C��L<K߅��8���Y�����HW׀�m�T<?{�2x'��k�}�p,��Sz����/���g6/ 6$�9���]Ш	����6� ���1C6�2��`���d�U�y7�䦄p�bUTS� lSۍ2�2Ͻ�X|f� H<O�)�A���e�3!d~ Wn��x
��Ͳ�	l*��+��� ���b u��;]~?ۍ�z��ӊ��4w���VN��I��{�[e�S!�f�/��H�)j-����!���\m�����M��S��5�$�:<�{K>H8�7m|Z~ht a�fq��s��߸����h����i�y���D����N�5o��;�l���m� }Di��(dq���O�)5�����di�a��Gx��㮭��=��5��Ϊ�\+�A~��_']s�0'SX��;4��'ba�x+|�*SZ�1?�����y�Ӷ�U����Ie���T�M�)h'�ʚ)'H�HI��E��_����3��f���ږL���~:l-3��Z~j����,����S�Dإ����p��/�t���6�����O�D?��tV�������\Ց:�ݟ�6(���O���G���g��=����*�S@/���̰b7Ӄ��إ�O��iq�����&�a�O&h� B��L�z�ӿ�9<�N���Y�ޚQ�S2�+7����f��D���7��Ng�e��C%ݫacz��Ky)A�FXH���:�\|����XD�I9���k���D�l���	Ʊ�������˴��Q�&*:��N0 �mUԛ��V�LZ�[P�@d�Ӑz���!���+�>��WhN�JuyV۸��Q�@@%V�.Z�l�ƃᕧ�E~E�J�T�2��jn�UoE���G!rB���s�Vȶ���ҀM�=bւ"��)Є]Mi=��酢˶'R���O��ո�e�l�]|''Ll�n5r9��q�bS4��aa��2c3�|��lX�ߢ{���4�.h�#|
�g,C��.�Ю!Ȟ��E)�t�}>�V�pX\k0δy}Gj�\����f��ZR�i3>��Z�3�9z��4b��AC�9�DW�Go|I:oP�種�6]l�*P�����C��A�k��I��a^���Yh��Fv��x%!iҙ��ݧ��4�Z�s�|94z�T�=��	����wD/.ѿ5��T(�"hh�/AC`b��o�i�������-�;��˖�w� h0eo'�VؙX���S,t#��*A&9 u4gv����!���v�a8N,W ��X�
����[�O�y�#̣+�d�K���X��$�x?ô�Q4�l����yY��+���¿P9��݁#��~5Zї�t�H�b�q�b��#m!��2��Z�i|�h�����a�ךּ���O�Tek}߀?v�K� ���PV$�6K&�R�9���*�����x߷�v�}ov��p���y<X���b��m�����?y�ͯ�4�D)����9<���q ���sF���|���'�5SS�ɠ�H9o�.��m�I�b(b�Y'��]�Q�Vyl:ړ�H�;e�����'jlh7�vd�J�]�X�nn��ܢ#�Q0s0qNЋ�38�07�~L�J����}0�kݏhj�[�m_�O?P�}-1�`�����
Xpk�$]?&e�#�[�F�����YU��|N[�4=o�:�)�a��2�~W~�e�����ȓlF��2᩟�Z�;��ɵ�Ivtg;�+��xjx�g!v�w�����sw KMp��������u�0P} �}�gX���s�"�B�p>c�����W��i��B�j�J�P�	���M�h`?���~�o�-���s�I=��}>�ü�=���5��>�r�0�@������f̗���C��|�6�"`���%��sR��I�QZh������ī^��g"\_?;|�;����ㇻ4�����p�UA�(�gf���m�?��aI���#Ҕ���=̷"9�Óa ;��"D�M��\�r��4��v�1�I����&EJ�L� y���Q�E��hOqt|�	r3$�Svg����Oᱸא� �Θ��%��u8v�].�p��]H��"E~���F:Έ�p���x:<�X�������F�q@��J�11R,Wy>�W��o���̄�^ �ך� 4Z�bP�Lq�)�hLV�H�!��� nĮE�CZ��Y1���7�3J����G�_�gc[4�����_X'���d?��sr���'�Np�-�۪-���s�zm���@U��mE/��dd��/���s���`��=�m��OUM��E�=�	9[R���i��ԫ���t:C���_Z�O���ѣ���H���mb�KT�2��n��*��3J�;?�h�Չ�zpI4���a����{���S3��ؗ�
��9̧A�_�)��>�|�\(��6�Q�e����Ty>�w�S�b9�,b!��K�Yr�H�׵\���˅�^���g�n����TPq�:�6+�(�R��x��I仼ʳ��YJ�l��BT>��W.f;e�	�����Jk�Pj�u����p�������S���/���j����Cy��vI���U��泭���$[�eFv0y�4| ��h��#�FO-ۦ�q&���ZX�H��Wd&a��
���$�
&5����:A�[��T���N2i���r�Nu�f	�$O�	��IZ<��|��x�o��ib<�E����� v������fw��3���Fn�����E-$���Zω���t%���Ѩ�&vo[r�n$���gXh	e�y�m�7��j!\�kpnr�{<ɚ�)0���8��v2�^9�T�"ԇ�ӵ��A4d���H?�bQ
�a}aq\T���@.�����D��R���,y�'w�K�!�9�b�aVw�e+�lIp2��%���#��`�˞�,q�i)�u}�>Nw-����Ij�^��&�X�P��bkZ�x�s��'+�g�ھ��@�'D�$s$��h�)ڄ-�5�'ߪ%��_i���$@d����Q�h�΂�8��ap,�L�I�C63G�(�a��n~�����^{a���ʃ���/�`��d��o0�%��=��O�L�I��C�㙕x�W`㑪�K���Jo�%�!iA*v{}�1���Ē
���!��t�-�Ug(�$�:Z�.Y[�0(0�����l�@��X>_Tѩ�����������
hD���^���+w��P<(]�����G�.'��U��,s �v"vb\�K�	
�X�X-q�꛿Ƴ�6$�w��:��cV
~���N,R�/G��,�G'��[-��\*�u��;�I�Xp���)
��9ػV���e~�_��:�Q���&̵�;I:Y�^��{��gy�ޫ��a�A�U�S�^�;3D��l�BI�B�J��������}ר���-�0��kp��;71Ўzc�����ƙv\�H�RV4
{Z>m9�B�Ŭ��;���|@�J�Pe�#��'�������xAڨ���3;K$Y-�Ұ�i�ϞH���Æ�hV�ł�	�H��Q}]EO���Rb�l����>p$���<ѥ++�F�X��*�9�G���S:���6���9ʤ���l]�@@�0�ޡ:V��d��&Ƌ�
�,����ixE59�Q�I�w�=Ԫ�^>�T���7'�^�[��=/���6Ɨd�����sF�Vo�J�%	��j�:pw��Ǘ���YqC��a4���>Z�R>��t!Vp]�̮K���u�P#�!k�������<��#tcw������wü����&��-����!S�!�6����T�x;���~F��@P!�F̬��J@��H0�ef�X�X�Z�R~�6�ig2�Ƴ�I�~~�e �8��j%��y�&&�7�3c����}�,
�!�ME�� J��2���b���@%cp�d��L�}��A�5F������mf�I� 7+X��z#��7��)����Ŝ���]$ɧa��h,n��
���D�-v�!i�X�bq���d�	?I��:a7ҏ��#<ix��^���� ���њټ��u$�=��+��1
�Lb�|�"=�I�ǕnaU4���5n�Vn�ɓ)Rc���aa�C�w��ڥ��P�^��Y�g`��#�W4�z��$��t��޼{��U�ȁV�&gP��ؤ�@�
�?�e��gt�",�y���QA�Z1f�b��*�Ш���ZO�K&,����zE�]/����������4w8"͈eօ�a���f���(݌���ƕY�<u<Z��$]jW�f8�؁��C�u~^/�� �5>.��l�YM�'��e-K�:.w����' PKE��%3FT��rH%pl�B#d�m� �k��v����y<��
x�ݜF�K�!���퉛pw��ɔ�N�>bk�.�kL���P�=�M|�iŃ��i�ε��#��X��s��>/3=34������ߪ��eG�"r#�U(���O��iU�;��A:/\���)�ܿ1��x4~2Hָ�muB���";�F^Cs�W�D�%hp�B݁������ڤa�6[��iHN�o�us�Yڹ�T<�e&���׈+օ�M�|&�,��T���.�[��ݶ�.ѽ���:�>�ٝ�$�
`�0�]�P���K{�� ���j��,�����s�<�n�9h7B&�����֍a��ʷC(cAnP�z�ÎA�v����Aj�j����`֦f(u�dr����> �<Uq���Z���vPN}���ߩa�F�CN������jM[��F�래h(	֒�U��$����(��+L�,s �+	~SI傠�?
,��o��p>6�[���֌�p�R>x �PȬ���ݞɂ�ŲM��5(L3t'����E����WG7>�z>��;�
���s��@ux��:����J�O�J��1j�����P����@V�&Gv��?�ӀMV׆,j�I��d�1>A�u�<u�{��.��h�F��������8>F����m���+^����K�` �^�%���{$�Fc�xp�-�v ���"1Z3#�L�pI�;����o�p�X�Ջ�X�*��~����tq��3X�Y^2��Y�5T��4�����E��	�Xڞ�h�l�<��T�.�_�>��%W/�e#sH+#BcS�#���=]j�q����,zn��Gg{9UIb�gN(֤���犻�i�\?oи�/�J��2�:��O�=��3��Áw��Yr�j�-��N�s��"^M��jSu�lR�����8�ĲI�������`?(O �ٮ*S����=4��q�B܆.� (ޏz\���C�&��7A�[�QS�[Bj���L~��u�#b�_+DD{�si�}q����%��\��l�-�l�ۂ��Y�h�JF9����.7H��N�4��v�g�A���֢Nb�I�n��r`��>(�%�~�mz��a8Ƀ�����Ȃ�B	E���}A���CNz>tU�K"Ǖ>~�tJq����	��M�-��7�A=�����;���[0W�̘j_7�n�8��ue�k�^�ʤ8�u6A�6�o�I���y�N7��6��@RAד2w���Ɵ�^��ח���v;�d��)9c72/��_�J;$M�E��-_�G{4z�����&�F9��^�_0C�Ot���"�%j�N;����Oʚm�(�XT]�Kd�<��l� z�:Y �`8�I��-��x~5����*��&�mz���7��ֺ��д�s�df�`�56e��o���Ke��ܝ��fP���ꨌ��U�y�栏�Uc������m3��I�h��6���;����6�+��=A �����E�ZdD	MP�_�[�|��/<,�����v�\����8��9�Hz¡��*�?s����>[�?B�N^��lN2�$!A
f$����X8ݾ@�0���|����U-m�%�j��l�_ ��I��8�����χ8����N@VbƙP�+�:�R��5�D#�����D�`��ߤe�=�bK\�s��VB(�_K0��~��4-1܏�EF��~�/1���A�8"��-ꕳg�}�&�`�?�oK��z�xb��+4%yl��%Q<3n���P�.�^ik���̷x�6@�S�_ק���:�?߇�f�TA���"�TK�:O�`ݩh5��+Yk�@�3I	C����]ak(&�5��o�j2����.,Hf\�ԥ7��}(�v���4��bw�RN:0�-���Mԯ����aژ.�T���2.p��6-�ػdm"d��wX��{�"���bЬ�=Ht��wy�A�SL���ĸ�Q�ϐ�h�9	V4E�4D�� ��w�8BL��{y=��0P{�2T�X��-� `����w�aP��0��\�Hp��@x�`&��
ˤh��n�8���S���6�xT�A�sY�����Q��z�[��Z��2bK�S�Z�N*������*�} ̝������>J�|/}a��+�/�8k^��¼��^�9�'`���DE�]���~ռ|\E��l��i0�
�b*a�Z$��_�Y����}aw�BR��wKPn��v"֧	f#�ג����K$Tn�[�4�$[�/�&[
<R�}\"���rf���������%�C''/�8�E+��K(�i���4�ĸ:^�	k4���7K#ɖ�i�����M�w�8UO���w��7O�������՜~3����#�8Λ�4w^fN�����9>�E�Ca��dҔ�E�E�V������I�\��W(2�/��F���X�f��f�����*���c�eI7��ע��7��v=�$^BjQ�6��>t&�n>$Zb�����zS���Om3�J�lC��c���%�ȹm e�󼲸�r~��8��W�(]�)7����b�C��Y�^r
z