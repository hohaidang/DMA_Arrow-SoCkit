��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW������r�c�v�e�������Q�6�E��>��P�&�?6(���I�٠b�A���V��0f���;���i�c��\� ޣY>H�E��3Բ�W�S��Ÿ��Ǟ�H� �a�C��|�� �P�Y�v��K��b��g�?��w� 1)��9Қ9��}I,�/{����OF#(�����\x�XCמ'�è+C��4L�6
�e6�"�}�y�!�e��)��ܨ0�E;��]Q�rqR9ڥß� �#�	\�,&�$�XgLx�6J�D�L� 2�F�sό����4ԘLTCo=��'Q}����;q��A���0=de�� �:+®��[sY��l=��D��MAt�7Σ���=e�F0P���eԲE~0���ODB4=�?�?���}T�i����0�@$V��i3�ܛ[���גw:#��q(>;�X��hM�ѓ�#��P�I���b'��.SЇ�lؕ�\�<3\�L�6�٩��_?� ;�/8wޛ��?��@��	s>���8y�v����z/W�SV�`��w�	���Н���Uޑw�Tׁ��7�x�{�b4�ܗ�\�\�p�h1��]/b�ԯ�Ϭmg�$l�!���J�3��ԏ�t.��/���3��%��WZ���	O\�1 i�Ǣb���Y��W����6�����n��_���\�D�N�ΖZ��
����j�3M��U��\��I��/p[b��G�32�u\@��t=<H�^|�E�]�tMD�r[W{�Y%��ש��nڽ:9X���̡fE�ܙ�|�d<�r|�2g
#[0�wˈ�WP�	?(��T�o�l���w��1B���GK����輅A�v\r"ʜ�gW���w*ok�gj�V[Pl�,C5��� ��k�����KI��G6G4E�Jp��m�/��q�� �^~۟���x!�az+�������m��/�X�tM��TP^f��͛����BH�#�-�#R�`�^�sWLl�lر0֛�Ҩ��<+�%[Ǿ��$��,���X��ۅ���5�֡�Ql��e[m���Ri�2/��$x�J�/#��M`����l�h�N�
F���8�i���xO�lL�
)X�M���(�JU=V�j|�)����6*2�H����s�@��/�����t���X13D���[���Nsl
h;H��d���S
U�
��@W�?F�\�_ew�^KE�s�(Uv9W
y� �.�mS?T.�����-�)�`Ap�j0��ÍA�H��Y{J��$���4�l��n�(�&�WYI�T���bH9��ۂV��s�rO��&U�,�p�B;�޺�@>��̬[|�;�esPW��9`t�xP����က�{��M�?CS�D��P�O���s�������|~&�bܿk⟁����%.�d"�S2��| @��#��^3�(Iw�6q.Z��j���Zք'��2qR�#��17ɫ�Ng�z�60�Ihτ+?�n�8������7�)g��E�W�����9���<~��%����-[�ǌ����Wr�Ԃ�ې4<���EwD�� ?3�#\ C��QBz2<�{ӻ��!mk���w� �K3oI��o;��ʀ�������$�C}q�}��zd�����]�՞���I�`�
,�B���?Q��5b�M�b؅�H�����?6��QI{i�0�=i�Bj��	�Mpj�´���M�_�B��}d*����!��M�-���2�tnk�% �S�I��>
Q�)��<ܫW3>�N������C~��C��D62=jK2��Vk��[4+T�����������0)��y��p�)H_ⅳn�����P O5���4~�Y��HO�y/а~wx�>����8,a"@J�$�dYa�U���nZ���]��	��1���vQK,6Y���X[#����0�%��P��r3��	�S�`���A
>E|��?)��/���bV"s5�]vv�J�W�_�#��l�2�Zœ���⺶��H� RL.�G�B�P�q�Q �տVbLH��Mc������&V�!�4 Ap���9�uG��B�k���������RM.I8ZL��Q�}���O��0	H�;�Ƒ�6���dRTv��e��#Z���.�j��o����E��횙�� �M�v��z�*����e���c|��0kDWkGu���K��G�8���;��SXa�uƱ�m��]�*�v���8`yw)8��L���x,�`|�v���6��q�h㤞��(m��0�>�"����݈�������:���X���h-X�@afнϴp Up��<�5����\eM���n�b�'t6����]	�z���3DDe��L�DN�өwTk�*��_�[JHp�=���G�#0?C��d��2{��vІ���s�A�^��3*ؿ���[GrĲ=��|��<�~ױ�<|����al�C�8�0ܯ.ͬvײc��_:�����Ф����+�}�IY��rqfUݵ���bb�C��mCh�7�;��/�?.�몺� ���05�L���i���� C��%�մ@�YB}�!$���TVx+^l䙁Hz����Q`xA\�>�	.s(�c*\���U ˲܅5�W�X������n�S8���m� <a������u�x�bp
�{�!�Wq�fWM�����Ŕ��&�B-�<2�f�.�R����a?����N�'} �VSC���7�)��o��&_�������[���J~��o�P��P4���=f|
0� jqE]�3�}�uD�Y��ה?E�����z/��B
�O
ѧ\YB�������0A���T�ǡF�ƹN�|n��[*���.�a?2�`X�;�p�tܶ��˾��@s��c���@]}q3�ܽ~B�5O�J�_8|��a���Ed�v�#�z,���"��o*٠m�LFa7�K'ۤ�+6�S���3t`٢@ɻG6"�2�m�h[�e(�)/D�B��8&��2C�m���Z���%�ZnH�+�S�`�.��vP^{��B�ۮ�X�?���N4��⌵ma��&ķ��î�uRKȲ��i��?�Xw�fu��]i'�h���]�w��X�tQ��Sd�U�lT"�v�cQ��$~�r/k,4��/~<��p@� �G�4���n5�t�� w9�Z�860��cSh�Ҵ�4^Ң��}_�ט�Cɳ��(��c�I��S7;N�5��+��6��&6_4���&�;˯[cۺ�5�󼾆���7tLI�U�hx��Hݏ�@���J{�0=��= 6�x7��}QM5��>!�W�E��1{�6�/@��H�N⤗��8��6�|g�����o��ֹM^�����Ƽ�zCbFv����G��*'-̤C�uA��{����Q�<���|�?H����0Q��Ы��Iv��̛�D�c�Ǭ�Ev�tg�>4c�p��G�p=�+��su�@��+6�ł�($_R$K�d���z&tXk惕���p֬O�ֶq��r�*�
�P��R�>���ꪭ�m�Dܬ����m��5��J�z%��εc�xh��
+L����gp���6�p���r��#���.΀Cvg
�҇Q@�t����EG2�Q�.��������pN$���i�^h\jt�[?�O�XED�݉Si��T�C��b97QI��~0rԕ!A�BS�_CZ���~��R룋�]��p����䅗ei����Gvh�8�%4�I�����x��0UO�}w	(i����	��,���@����zy��&4��;:�TY�iT�^e�*�ӯE�Y�$��\94P�.�G0h
��.���L^r��E�M�}'w[1��$�ݫ��|iq5efa�����&�g����idBbd9{�u�]��Hy�DL���z����m�Q���j�ŴU�H��p�rM~v�p3�$Ÿj�8�����[�\����%��4 �q!wU.9�\kP�.��%x?��c�氣�>�gBG����-��%�2W.��y�q�"M���5���f-�J��% 	E^f�յ��_�Y��;��;p�*�./���۟XT���4�6򳫡l�X7S�I���z^�Loг�����^�&h��q[���,�}!x�!\�2�L#���kR����3}$�x�#.�K�vE���G8�ƌY|��rC������R0����}-�����lOR�#�cv��|�;����2_� ��<s���q��Ԅ�K��x�=D�lW2��;F���ёƌ�B��]�:D`�'T7���N�i���IrX�	�@�b�6��m��.ߘ+�[�B��[����CCIY?&���$�m=q�
!�Xzxa���W��� �X5�9缗ɝRF�L�?Z�H|�'���q҂��U9�{�|�M���H{sD�Xūp���D"B�8n�V�Mn�,蝡<��S��DI�v���Vc�_�;���^~
A�0���q�N�������Dɕ��.���|I?Pm���A�	�@�;V�е��+��6f�l���k
4�q@qL�V�VJ��]&���z�n�֦�m!�'e�)q�M)�{�`;�:/��s�S8Vz���1�m����o�"mǗQ������I%�vצh�^�Fz������RiZ6���Υ�x�J�l�=��6� LnFİ�a�^&M�I�P"@���_��S�b
�k�bz(��%�0X�J7�������ගJϦ8����A�q�:�0��
�`U��h��ڿ���F����l��	��˂z~I����)��$��k
6#��A�z"�YΣ+�>���;��C���c��l��4
��h�$300< �8��C%$�~b�Wi����B��f�t�����̖b��<��쁵�s���NSiQ�X(������c}'X3��A:aނגH�ެQ�7ݏ@���r#�vVGqF@Y��Ǻ9	M�f�{'^������wl"��=��HO\�PGh:�,���Y�ag"r�_��-�kC���2��T=�[��[��Y�R�PpE�_�L��L�W�4�O-�H��)�`2(�OP$yt3 ��;���>��Y@w=�Kb�<���d�[���B\��4���N�o������bQ����B�}�B���}��z4��2�q�}���c�<Vǟ�4}�7'�!z�N��A��b�1��\�0�H�6�O���:�0�߱g{;�/lx�KV��ńan�^�p����b���i��b�f�cp�yqf���G��I����>�2��"���e	���v5J�sd�z^�N8z��_�"OK��)�����r�3���}ÃjK6�=C�h`L��Nޠ\j��#�͠{��u��I;� {��9���	0�n�ͨ�r�����_ʕ�5�{TM���*d� 	JU��b?-q�^H��;P�՞�ay,lJD:

��0ncƢ������Cʼ[;����Gi�|L�Q����W�L���j�����}�=�;?�l$�Igj�<�}	��a��j�5���<������:XP�N&>�9���)"S���.1҇�i��Aմ��~E��a�����L��=E�Q,QB������8�X�����x8'S.b��l�i���{����xNh�y�Zǻ��y�׾�\&��obeN��P�uYB��9z��!�eX��z[H�
T��Dv_�ٓ쩀0w#��|)FX���ĜZ���.�a�W��I�������hj��*wM���}�3w}��֫���U�Z�ũ���E��5`�tp�E���d׊��{%�mf�ϕdظrWwp�Ґ��� #��l^�|Cqg?�3|�Y�M׊�kr�KAw]�-�Sg��_y"[�٨c��)�wM�}JDh��#s������	��_Q,왬�/<��;�Yj��rԯ~mRm^���R˿>�|ݤP�|�M����C�$8((��r�=�	te�&D���aRI�*��?��[�!�&/�;����O^7S&�>W���
����sV��*5���EG\`�td6�_ɖ����H9 �q�p5K}Qk/CM���Z�xJ���E'GH����<*uҧ	H�)hK��ګ�m=��@۹e��H/�3UE��#���i�w>�+����9������s�Q{>X�Ur�I��ީhۓz�{��潏_}��6�9��IضV���O�g�<�􎺃Iv���J���|o`z��e.瑞-�׏�p��=nݯ!ʜ&�ս6��O�<���X�
e�0���J�0�����Av���|�D%���|��P��%��T�p��j�s��6���A��H�s��_ō�]aS�����FDQj�i [>"��sT�o:?T�5b�l���f���?'E�{��K��rDs�U�c��c�	Yu�#YP�
 'o�w3v��f���6���x=�$M�l�t��9\�Úr"�n(�F�>�:��j�[^|n�K�6��1��{;>����r�}cf1�ݞ:�ߒ �pY�5����9"��56��g�+�54��!�&����D�������<�h ��D
�N+ ��L��ZƘ����'����1K�\iݕ�<D��$#m��7P[��?JJo��P�+�{�q�}��F��H�A����p��e�-�3С��f�U�щ�?����od�(��grB,���J1@4����-���/j`�T@N>��W��R�;,!�h����9��8DU|'��ܶ��9�L�qqJ �CV��T������ӋO�Z�fͭ���)�v,��Z��#�C��ǈճ���3Lm���j�=����Q��g� �O��4����m_�.����)��t,�E��2����s����Z�y𬈣�.gq�CyB��ϴt����K��-,9F�Ϝ�d�b��7�/�"��znN��+�F�B�a�z��g7�A�
�q[��	/κy����ٯ�*#VhʭG'�������x��'W�=A�E���b�����E�� ����y#x�d���(�޴ٚ<(*��- �s���=#ܼ��7-燺�K;��,q(.��  �ɺj������=��Z�B���n�jA��\�F�1Xgqň���F�s���K�>��Zפp�<f6��*#�4JV��>3#�	�ރo��뤻
Ѥ�Q5�r;gl�A	���~����y�F�U�>+�����[P06��r�����-T-h�E,�v5ܕ�]��h>���ѭ�!�=��`���D�[4�`"�L����|�f8�߹�U��n3��2��tˀ5��ըb�P�nK�]�����K����e+��|nO�j�2��"�\fץV�M�=Mh��н�Y�g�N \�э���o��8n�]j��Y$:�ogH�\,�z1.����0��/^��c#���!dɃ2+"���J��ڢ�)�ƹ9�@&�:���>�0�Q�xK^���؞�����@��Nv��N���JM�6uQ~H�����=�sk73vo���(����G�'�_�k�2��� ���q�kΦZ�5�Gt#�W���O����'Ǆ� Ip�7Z6�2���XN]���\v�?�R>�v-MU�'�� 	��s�u��LI�{(��Q"~&.װV?�����=�>�=NV�� ܚ?�b�B\����ЮW>�X��ʌ������'��?���R�}����&��q��K���C�j�8d`��t�!����&X;�br�����7�B���̣��T���wvNp��݅ʑ�9��u0��\wܾ�XJ�5ĵ>Tzh��e��4:+vY�5�O��zp�l���}�3�K
���H��@;�u9�����K�\�f���N��:�I���X���J�v�aE��|%>T��aAtX��@�L���8(Hhb��?'~������o/~/�<�^�ۀ9O��m����C�dg���Y]sT��]�٣�b�x=��A)h��o����NO�D���Ԃ�r\�
EKխ��[2u��LSU9�z!��mG^�\�g|=X���RTpJ���ZHS��lw؛2م��q#����AfV�df��,�ݪݰ#�S2��O���$F���6Ƭl���,>� >�v?Z��a*�D47s��'��C˰�Z�d��l��3��p��	^ˆ?�T�<NLW���� }!��N��5<D�S��j������_�_e���\�.�]N��3�t�5#vj�����cmG�)&$��/�C��LwB��/6�C��˃���n/LkǴ�gHQ"�-1�����I�v ;
��B��:�9��;.�p�_@��ڀ�Q��?�E�KĖ�3ү*��Bve�Y�Ä�O{��DtD@3�RZC���>3!�QoTy�֜�n+%�����yC��?^�gżIz��DǜGMa��e'r�j�c��5S$qh��C��حIh
������ �=1l��Y��LG������cf3E"=��W�:��F���fv銔������ȟ�3t{zD}����#_N���x7��B*�a�o�����$�m�����@�+��V�of(�����;�@�����
I�h
[Ey��t�uh�Mr�����f������.�qpM!7�"��Q��Mx��2�2 j�k�Ɍ���>�UmJ ;�H=�_gY��W�W���%�4a�_��|Yt�>O4�1W
�ą�ObC9�筬��5Wk$d�*}q1���(y*:�M'�2�<F��3�uQ��?@������`��ͬ_��������D�
͕c��t������"�|���϶+JOGK��J
X�]w&�N|��+.�8Sa�~�:�˛��M@v��\5��Q p|<�Lj���ƨ?�w��\]x����(�H��5�7.n,ac!�ݍ��3t7=�\-"v��H�=u{���t!Yq��ZA��p �}R�J�		T� ��]�V�_k<ՙ�5��!c\�F�F��)r�������W�G�k�K�(^Y���S��J��ȫ����z)�s]�gu}7I�eBV[zX2�t����=��Q(r��ߥ/X�u�V�����t��'�������iZ��c�&խͅ�QIZB����
��;~{���A���{��"G_?��������-�>CÙ�$$�1��N��5t�8ℤ��uu+����X��#� ]o�1�!�Nz����A �pt��Q���o	��=]
?�ӮJo�ʡ��a����O,����t'~C!��<q�f�FR������ظi(�'?>n�J��g��a	�#J|�!�RXnm8��=�������v���D�߰��"����I6q��:����K)o����y��i�%2����b�9��&���������I*��c�!w�kMd��*0��H�i�/���چZ�F��<�|��IpQU�Q*��ڡ�� �c8' Y�2w[6
p�`a�L��brCRE��F�1�������� �ȁ��i+:5+V�5�Y;��`��l��P3=������$�4q:��4΁���E
ư@���M���63�� ������Et:��g&�b����C`i���L�6�D �$��9Fܚ/\�L�K��f[���g��)ւɜ��;T��'۪ߛSO��k��|�;���M5���5U5�uq3��d�����ƻQYm�5����oc�|W+l��ٵU�	V��O���5dy�&,;�=-���-���ZE"D>D��%�m�i3�����GF�n^�Qs���6���^Y�F̢��Hn��V�>������w�O�-��It���)T/�c7NxGe@�+��Be��:��)�+\ ���3�;�hփ#�KwJf�R�l��t߉� ���(ҥ>x��V!c��$V��>���j��Ѩǲ�*^΃�;�2���-3g�YN��H��=E��X�����4�	bURC�TY��H���E���h?d����5n?��f�����b�b�u�CE8Z�����q�����P�d�
U*��Kd��!K���Ji\��#1i�d%��T\�U����>�b���#i<ní����*������~�]LO�ao��n���уM�~�q�%r4j�2��Cv���'��(����x����_�O��E�z�a�����cֹcR�f0�"�8�tk��xa��ԥ � �mؔ�n� ��E��cG.G5���@����@$l����-7�1d��kDM0X��W�Ggu�ݬ���PP�kY�F�:�}��4E'D%����p����A�cj:L\h�K�^P��ZS����y� r���\�C��Z�ohrүq�V��H,QڭM|�jIK�z�����׉T�]N�Cc��q�Ey�z���c�уә"�u&�آ2r�0���Z����vN|n?�nrʤh{���-Ы��r�B��m��n��Rae���?�<�q�ס�ԙ~�9*��7|K˿�G�Ģ+���<4�J���ji��PB�,�F�Ձp��?.�}�w֎5�o|F����ƼƿQ��Uv@.��`�q������%K�~cd���f�����6� �ҼXm����Kƃ2�pe�Ü?s�JW���|B��=�6m���ߕw�j{5���dV�,�|�61᥊�Sg�k��`_�c�� �g���
R���B�����@!$�h�$��������4�]4r��o�˳z�Է�o��;��})HW�ŭh� a\�B/�	�n�q��'�Q�hI'Ha�e�Ŋ��Qaֶs�M���z��_�Xp0���]���8Q@,y�U���ëW����D��+Z�_CM��t��qa���j���{t��I����<����_J����-�_М�#��o��/�5��8�6����׎��+qk�ں���?�Y|���YA�k��}���*�1A�� ȓ�����I�Gw�a�a�Z_*[֩�s�Z�j ��д��a0��T�(���DY`����ݱ�
��Ͼ������&Ek@��R�J5�+����s�P1�
��/+'�=� ���Gt�2fM����p�͇`ؕ��N�4�:��$̬!���?��&åL�� 6�̌� J��v�u�m � ;]�NE��E�@t��� �$z-kRR�pC�-1�%�v!�n2K��gO�13�>�<9�d鑤�Ä�I޶���	�7�K�ۗS4��tre���(�A_p	�wɘv(|k������9?C��C���y^2L�g�w90Q����g�a��:a�����d�aw#�i)� 4�(k-l�n̕=K�2�lO6�dUk ����N�i(�����á�Q���a�U	�9��&����C�s$���uH؏�v��yP�G��(��9-z#R-���x�7��%A(�D.�sl�t�zI�����($+���i�6[�T%�@��}��/�{�ul�g{��D����_GX��:���F�5��zU��Zh�e���&�Y��8���d>74�^���ِ;L�b<>���,	~�x�L�'su��.�њ����Y� ���q�{:�^��L������_��+%Ƈ�)E>�Y�#��u��\@�x����j���@�|��Ħ��a�ß�v��4�����v
����t�}·�>U�����rd�tn���D3��s��ԉ)�	��߶��.�����X�F��M�ZN���e֖�4��t��������s���/��?�L�����[�K|5�1�bv����t�.p���̋��з�I��zK7"�'͸O���|b�;<L�c�D���\�����"���^��J�+�ޞE�)�� �A_H7�cs!�7PV.����P�<��/$3�lڏ�{B�~3��<�tTb��P.�Bh)7\%�.5h��w��9����A��mz��Y�Fߜd7��pPӽ��[N��%�oN�.QӋ�
�� �諈�NZ�6�A�{'��D/��$�#�i�~h�8xV������4zG���,6�F�ѽ/���9��P���I��K�]T�偅iv����Ǝ���ݰ"Js��C�a�N��X��f�CE?|����]�����`���I�3�_�Z3�6�M���6Ǿ�l����v<6��}tA��h4g�c���>vM� ����>��O����;	��V�T���#2�ur��{�E����������#�v���.˥.D�a%|�O�;˄ ���%|f.n}�Q	Hλz�Y��+��*7ǝ/���dѿfd�Ԕw�Qoa�'~EBE�g/�_e�zn��ǿs͕l�M�P&���=�8���d�t3�T�Р����XɅ���O���H[�j����J�ӻ��QPÈ�M�4�cY���Cz������d$���hְ�[�c�)gF��L����To����4h�v�ag8�2}R�w7���za��?����ݦ't�U
z!������w�^���6o+)�'c��*��#+1�C�o�C)��
I�O����zo�]t���������$w�87C��T�a��WG>q�S̓|�s%mL�Ҵ��N�`p��/' g���
��=��T�T~�v�ֺ�z��Kb��z�@]qU�i�2�-l%�[)��a㛉�F�U�2O��0Fi��$%	5W ~��Oë��3YL ؉%W���:�!?�����Q��o,�.�uٹ�
Eƥ����3J�!�i��%�{��<�`ŋ[[I!$��W�-*�]�"���	�����a~�
��$��)�F����ˣq��i���H�Qw����S��6��%L�߃���n��љ�	�]�7�ه�������F�Ú!�ִ����TQ`��tn�㙀O����)IíFD�k-���W��U���N��jg:����54���ݵt�R�1��SBBm��z"��P�֝T�ݒ ot���2N[g1Qo�е/J�_�Kfp\�V�f�°��ԗ̀�sS:]�\�26PS���P�1b�[|-xc��Pw�n�d=v��uVﾌ�Q����N-=�6;��*�C-;8�Pm憰
�v�#��z��+���[��8���9��=�_�u��1��x>7��QQ���jԫ&nD�`h��2��J��']�����O�N1je�t(:Q2SJD�^�e�*U�.��}s��!b)��_b
��Fe%�q��usIW��x�8<C�Bm���ΜD:��l	�ϛ��֨���B_e�h��Y��$tz���F~8m]j�������z13�M�\��*��5��*������=��P���#x]Q �3�Q`տ�d�9��t7�~w8c��O�f���P��g�O7�q������e���,и���\ �G�O��s��,d�BWH-v§}QC-�4�*	�y	Uqt̆o3J/3�q"Gw�����oY25S�Ҳ�֋�v*��;���p��N�S����k��g��42�!(a1�i��K�^��W~j[vո����}������� �wzjڷ�!����N�$)/���B�C���q0�ѕds�!ht[rO,���`�=:^@�v	�64=BrVAv��{�.�B;�v7�X�O�������^Z�tƾDD��PX�hD� �-򊀙f��o$�t{�mv��Q�rӰ*x��+��Rl\�0g����[mhS����Y%���fX�����;&�AU�+*K��F��\ϸ\lʾvx,��1b�2g��(\M�\z�?�2�	�	[i��=��q%�bD!���/�`Χ�KK�0x�Y���6x�Kr�z�au���ê=�p:�m�(u,D3�����Fs�Q��9� v�����os+Y���*��(y)���`\Dѣ��
`���U\?ãCZ��㎸��n3S�:����� �ݢ�tc���?�������{�٤�FTp�������$>�[�7�*8H6 �׈�FY��KHK�(9���Qz��_Ց@Sp�0��~a���c�XK�3a��feC-��J��ԍ+?B�\��WH��m�+Ų��e�N�,p^?K+��e�,�8�G�^�2�6����f�~��R�q�F�גz��&���V~�֮�9,C�����,�w�ON�9Ŧ<�j|�	@���D���������։��p�K71�K�"�;��")��'��[ |fs�f�~�EW�.0�^K!��Tǵ0�VWg)%gQ	�����5@�1 �јwo9V���{�~��#��9������0��
����k��L��=b�3����cZ�'8���š�jdP�/�|[�g��8>�T�����Ix�����.���j���Y��p�K,9\ֹV��p7z��G{�a����ڻ�4`��,�p-�m�j�cv@
Q-
i�j�)�
W����_U�I����e�P�;~�4󧼪"���pMo�(D�	�w����j���K
8�[��ֶӮ�R�h	�:I;;��m�4 �E��&2 q��-[8"��0�4��m$����D�����@u}�XJ���l�֖Y\�2A ��6@�ϝؗ|��|p�7�m�1�!���i�;O���=ǩ�(΃u��Wdz����̔�Z,^�l�F��B�6�_6�d\���5br�<�JKAD5�M�qvNu�x<b�h ��3��pe'�EP_� %f�/4v8)���;�h#wK�6w��6wFFR+�0�T�	�(iax*9�����~�w'

*J���M�"�*]5ns��Q��\Қȋ:��=�
/���P����DT+/E~wO��C��<^�~�\p�����K_��+X����趤Ao��P����%�1���X!Vq��^a�O1!�&�fRK@Z���:4�<��Ψ��"$jV����7K�̊�����������w�~8@�p�4ޮS{y	�Y�=�|.��ˑ������mp+*��I�䰪�d��Q�*���hȾf D����>�iKr)�Ǔ��������0�Lc�Kҵǩۦ�'�Kgmns��R:�\�#r y@,�>�j�X�qG� �����(h���^fNlϨ�� ���ǃ'W�R "�H9v3�VcӬ�B�v���6�}������R@C�{��;����;+
"�r�s`��F�Tj
M��n�m=�W>���k'nk���p��<�� �>U�����x�e8v
����!�uJ�0P�6�����uy�{����z�~�W��G�����%A����^��j2/I˃�r(E�t���/��m�`͐p�#�X���P�����g����-�1΂EDDe�N��G�����#a-z��"o�YY@`����$�~J�`��X{߷YE�D��4/��Z�ti���кS#�P���:�N��B�6�%,��^�/%݃!�{�.@���/�Z�n��jM�`�Ĵ�.��d)��b�6P���(���Ҝ�׌��>T��UwO��{&T:�6�LF�v"�C��qQ�^�/�Cp����.K��\5��I��	G�8FA��rg��us�F������z:'����y_�ʠ͞_:�������KJ��{�CgLN���Z+)�16���<;^?�:����WYײ82��p���Q�4vT�,`�����(��խ�94J%8t��T�
���8����`�dH�lZ�� ��8)�IT��{Hm�>C~�A�v�n]_(f��Hj��AvW�ֹ�M�.^�B�' �|I�׹!13��)1b���eP�~}?R"U�e�#j�Mع}r�,P�������Oon�9�13ի+B+�����;��$D���S�J�;�it�����Wd8�x"������ ��$�tF[��=Fp|B�T�	vswTK������@��>�\bBԆ4w$���0Ã\	{7�,����L��Vl���55�Ow��/�Eo�x������ ��|����T��T"� i��������?�Z�R2:Ϫk1?sg�!�%d��T�rPՓ�|�x֋۔�q��=�y�r�F.����b��y�X״���s���B�j#��:N=���>��h��5���aw����/S9����� �ic��?�4@9\���,�N�j�7�l��~ʝ����0 !�t��-?�k�P2{rƸ@j*�&"�Ƕg`˓W9��mo���D�o���_B����*{r�=��0�]aТ�(���h�!D"8�C\N|�V�yꋽ�Ƙ�u"@Ҫ�����]���*ą����Xo���봃 K�~Y���ݸό��k�7�8:0a糃X�<_Wi��M��0��m���9.EH�~��	�ѭ��FA�OPp`�2����+D3/s� z�-���X�n��ά��6e�3h�p��ɠ$	����ң�6e#z�ȕ�J�k��x�t=S��p3E�%ْ���!��'�v����@�E.g�X�d	�*�8/Z��cV�w���d�������Fs�
��k��ZL��|�:��^e��,��GvM ɥhsV�V�n�Z)ћ����x��O�s'ĹS[~w���LB�x���̦\C�\e��}��$t~��0$O���n ��zsR4��b�
I ��'��g�����C��[��$�-&r�҄S<�i�Ug F��i�C��m�u��J����t���?��� ,#�T���mL sy��h�)�fQ��B r!�
��T]"XqͲc�x�R��������R�v4J�#rW��Đ޻�<ɉ�eG�}��z�F�Tw�5�Ȥ�h��������O�z���{�������k�_���@���>��y/_�}hQ�U�>��S�H�j˷����"�hz�Y�N�Dʱ��A�ې+��9Q�Ƨs�>��%��s�\�v�>|�xǯ$�l@b ��Y�b��@��̴@&z� Ƶ�G֊[���ȋO&�kd��90��Y����ܽ�c�+��w)Xh�ep@Xg7�O
��X�B�R�p�W�ʹ��Ն�I?���*y���^"�B�M?�q:�_���}P�C�?+nH�"#�����?�]Ah���p���j=K��mo�S�\]�@��C�Dh��B��q��r1� :Q�<Na�ж�ܸ?��$_Y�Ij�~���y�F�#�w�uf�%\Xz�µ���FТI`O�%qP3cJ����c�q�k!��E�ab�����)~���u�oH����d�8��� "�$��K�`�v��B�t�8�՛�=+��o�%O�x��W�F�P��篘��A� ��D�)�mݭᙎ�ҥL���±�U�������%N3�uat7_�!N�:�ć�_{֭H	�L;؈�)d��}�}:�WHpђ�f\*OiZ �������tбP#�4m�C��
�����s(�ȇ�/�8oG%�+ee.�9T�����(����1�Β�s<�����x�O�������v|{u����>q8�g�ۗ}u,e%z7�-�Go�=����� bt�TO�@�[�_-宪;"3?s�G�ކzW�ٙ[�L�H�n���Gk��sӈ-w.�����D�����#�_��F�W����E�h߇z�[E��Ct�hqN��ՙ�ޚe����o��
Fi�e�=w�U�u
rt+�xD�B��}���k�ψC�����x����3JwVe�u��r��ER��;+���Ar�S��'�l��$�5m�\�<����O.E<���|�%pn6r!!�;�c���V����ch������}�EDM����^&ڣ��L�'��(��(n�"�H�U�����嗀 @M��$#�pV�Ho��gE+-O6��+�N�Y#�%�Y1{�1��Y���{:]�CV-r�1Ɉ*N�K-�[*`K�5U���"����mDPmBT�/ʡ��Q�r��c6N��xM�x�3+Zg������qa�D������u���i���W@�Hx}Gt��7vV~w>��ԥ�1c��Gq�w���Y�(�i:�jPV=�uX�88������ kJ9�=�Cm�\A����yAŌ	���K�L�Dfه
ol����U�/P�05
O*s,L�߁Uy�W�V5�}Z�}C�w�&�ᾰ"����]Ǜ ��P��ܐ��&0�8�vB����	�fq�jdbױE�����&�����f�Sn K�Ӛԇ����P-۴SQ��wr��`	��\�l�%)��:�$�Rj�j�ğW��OٶF�`߿��+7��
`�xY�"���ܥ)+��N|I����Z�����6�dlR��^�b���`tX+٪���$Yf����ݵ���]S�y�!�^��X�y�Q��4�)�l���%ΨFt���l�R�̞w�1�p�\S����2�8n!>/�W�4�t�Z5��K�J^�͑�[�L6���̙��	�2KC3�=�w�#ĐD�(j)��N�{ѭ�h��1|o�_��\?�3�Oci���+$� #�!%c:�C.��KK�J���7t*JJ?QT�;��ޏ�!��ϠJQ��Ç�m l�Un�̩X�ѯ��PsߺT�utt9�ڱ?�b�Y�K�/P�wgh����Q�������'�g���#qx렿yi�Z��(�1�]G����6��L	���;�:�S��x�ʴm5��y�<��e5��7�׭���X8���u�W!���ang׈�0 j�l�_R{��h�� I�RC�H�p|�����Z���N�H�w�������͕��Zb��³s�Z�4W~�ϬIoq��:����"͂��@Ri��>+}4;��c�d2�3t�E���Z�e@A���	;��8�T��ܤ���6,-�k{�5�)OQ���K��=���/�����$�ܯ�����m��|
�X+�\��ւƼ��~��	�����z9Ewמ��Pt.�ت`U0�����+�\+��F�G���}
��c�G}%{��ӳ�|��@Y��e�_�AIi�/�ʧ��%��r���%�eU~��c&s>����z����2�M5���!��d�zxg]	�LX��"i�dy�:�!D� )��([l�sP1F���gT��k"����Ue�h��<D�$* ��:����zP�ⴇe���p�f�V�>ܥ+ ӓ!,}m��6���l�E�Dm��}��Ķ{�O钌�����"���'�+M���̮�i����2r��SV��
^g��Z�f|�#���~<[�=� �Q��!�Xl#��1�$~��P����������N`�q��zM-+��˳�x\���zŔ8�b��;�o�b�-KZ{Lj�Х����4�ٗ�k�0x��"�DI�d��]��xF��q��S^�=�&˿ݣ@������m����iԼ.�^�]���&,gX[�s	~-T�ƈ��`�pb'Q��� X�廋y�=���k�� �R���p�s����<{p��xGK��TG�w�j�	�c�e8Aә�F��x��y*a
�6��)fUlq^o�:�唓�M<��g�9У���l����������	��ʣ�;Ӎ��1��=�'�F��x�P��]ʦ��`w#;f`3C�TA���{R*>��z{�@�Is��h�z����/V�M�($@�� f��׿�b�l{�����В�K"m\�/������J�$<�S9�=|6�rZ�y9�u71��E�L���` )0����g���+j�+��X�ޯ��F��ҽ���w,+�HT���cm��wêr����9��m���-
+�����6���3E)-
3Dy�B��{�*-��̺�|�����`�GE"5r�zf@R�;
�T1й�����S�6r��bQ��IE��Z?�B[��-�|xT����.4].쨃o���h"��k~4L�ÓE/�K��s�>c	�ׁd������XR3���S�X-���C��Tj���F&��'լ��\�]a�r���aF�S�i�4u4ӡy��#늷NR��X}���v�4M�Vq��_`I�+�V�Q�$Fa�#�;��4c�ْv�W�*��o\68��������OEϴ�::@��?	]:�7!�H�@�-�pA|q�?P���]��t��_�����+û:Nn��7��C�̄�_~�2<��r��d�������� �a�}�=��*�K������ѐ��k�%�l�¿��(�C�
��P�{>=�U����'3?�$6�0"�����:Ѳţm�gO�݌�N�\��Ë.L��@�5��`��4��1�D�KM�O'�xFN��$�9h��i��%G�.:�
�L�@h]��90�����fC_�4�� �+(��gj�-'�%D b�*E��ob�[O+�ݧaxɶ�AL�e���ز ���:�G�{zy -�U�	FW&03�(��bJf��Uq@%f������/=��2$}���W�w�?����!_h��&��q���G�n�c2·>�-|q��Cy��-v���8h�>��~ ��1�;�K�Υ���n�z�+��ِmѨ˿���Ŀ�յ�X˾�G�{Y>���iygگbx��K9�-#�ofkY�¹5���&6J�C$�%���1OR����
�2nPK�HQ��gw�4aD��K�����6~�/����֌���r*Ŵ����Wu�Q�[*��#���Wmo����E$����kt�i��r�w���d�iK���J�7HL:�4�c�R�3lh�j���
��c�*�gx]�����}:-�UIj]z�F�u�7W�jSQ'��o����^य/�N^6���$E񘗯�|�W��Y{H�j_�4�e�_t�׸t�[��-��g(y��)�e��b��M��Χr�$N�9[=
��8�.9�*��P��%�6�C:l�q�T��bwr�0w�~���1ش�j����`�,����ko:���]���o�^0f؃c�9*Z�]+G���Xd�,���ya��6���f�T�2���lM@���L�͘xq�q��c������0�Y�����<�L����2�^�jZ�KuRpMȽ����x�)S�r8�a+�	�u�)(Ǎ��^]ASH2�}i�9��zA��~��@����*�2�.�k��e��}P��O̬��(.�O�Ze�c[�����ܟ�T����A�,�J`��w���4����ٙu�:P��x	�I����� K}�U���f�]a}40j�|��!���>��oǚ���>4����/�>�̼�L�������u*WBV�h{���]>@9+���O�cغ�1�[�ieEG\(��}eyI�ƿ2�� �9ԍf�� 
v�e���L'�d����$.�s=�4v����|\�g���p�Yh�iY�[�~N�o���D�ReY��.5�E�(f%J1��v�2&��49�n>4��`n@�gԹw��+��l�TK�d3��S;�E�K�A}���Ϧ��i��+�"O]�z:nԱ0��ʕ�m�#HAZz��܀e����$�b�Y�h�U�)>zb#��W��L�r���` p��z����^|���#/gP	h3��&x@<���*-����S"J����x�.
A
��s�qkZ����W��8b�\���Y�fc~��!��Y�b�Z��*������l/��s�ט��ےD��j�@Me��|�Pm�m����@���l�$&���Qg�O�><���
�nd��y����\�S�^(=��h�o�����k<�aϏ���)��#Xoa���� �-X����Ԟ;xvzZ��z
�u��@��3`�V9_��
>�1WЄ��1��/� �<� ����A�b4�*�}����ah�c��iH��n'��Su�y�����ju`v���\�AS<�p����vN�s]��_���{�[o�^���릖^���!��>H��P��lF���e�9�f_�gZ���	PScDz��$RWr0�;�p�;T	Kb]ۀ1��s�a|����K�gR�.��Y�C����	���I�~������ҫz���ʽ#��Η.��
��~>Q�A.5~�{��4�bm}u/��� ����pW�@t� '`��<���O#�!��7�u=O���l�������Cj�� -�9��t��]�q)d�> 4����|Xs�np�L��F��4}H�6통7:��c�Iy�>����댞
�s>e�����?Zv���:������,�O��K�I3BC�.�zҹo�,�!�ɶ�qߓ@2n�	����:�lM*ڞ���c\���<���=�Q�S�^���|�<�����#᭢Ȑl\�[Y4��8	G�lE���R�`�)�k�(sQG!���S�[5�\"����<򀪊+j"�"�=f��� ����ɰ`���߅�$h�ݧ��t@�r�`��|�L�\��w��HS�(����L����o����]P�C�h����du<�`3]u�m4X�5❩�$��3*F%���F���F��R:!��\�L����X�}������ü▢��� ��k��b@ǃ6�LC����w
��ޮ��1���INm��K\2����۟�Z���B��zG�؉o���Cթ��#�B޳��y;/�ٺǴ����U�H���}{��̪����~�0�b�G�R�nI���?���G�g8��"�y�����F3~�s�dx�]��h;�;��<%&�p���^�H����!�Z��+����M�S��|'�
��B�*#�!i�J�,�ڀRͨm�η$0uRm�v�m�i��`sz3h�V)��7X��4d�1���K����lZ]���i�"�S�*͓�a�w�S�����:y�~�Fd��O�;$�� ?�y݊�Ӧ��B��vA֨��l��8�d��l��8#��4������]QX��-_�o>��h�E���Z��ج�=%�F2�~06t̑�,;4%��m&��.��Uc{���v@"+bHo �0�}yFs{;h�8�B]��~_�.�O�Q�*?ܕ�<�<Ⱋ
܄���^��	����ا+ �Ṽ�!���}�G���ӂ�4HذO(o�U�j����������G&�T���(�����1PGK����<����ž���17YKugh���͆�waR�H{��y���`�*k;& �̄}���
q~����[	��7t���4�����2O|��R�R+#)΍U���%lEAF�=\s��Z3މ�cm�1|����A�ǹ)���Mq�:��b/x�y��P/��ic	(�%�v�i9X<����
�J����_0��{A3(�����ߔr��,q��}L;�8��S~�s�^�vQ2����AE����qҠB��:���ɐo�N��_Mo|vD���To���]��e6M���[AM�Ѳ��Uh�C����+X�	��$�~�E�M8�գI����C_u��_8A-���z���ދo�s�~��J��W��ټҚ@/�,z �J[_���Z$W(~�$@�`�{-~kѷ�b	��:�QKs�bDx3���GAt:pDtF�
�d#����4��3���W��cy����hH翮�b����%clٲ�x-'���UW!J��Yh���i�Ҷ�V���N&���ި$ �������vSRt�1��?(;�-��5�&6�L��ïFݘ�Z��o9��Dޥ&o|`L�33U�-f���W���A�YxX�W�8�8t�x��=KzN�k��)`M�3*1<�K�ش���~@p�9�	��(� ��qْ
��c�s���͗�������ǝg�I��O{�����>�S�D�":q]pf�&EGԻ���<���=����5r(s����=yO�h�j�h�؛yō�&�K�mS؇�g�3v���Ƣ�`G�t5NׁKO��Vsϱ^�ف�I�)P�m{�EMż���V�(�16����䫕�!�G�>�h��%A�.�='t; �Io5xy��&W��.�4��h��[\獿P1Pῷ�m���z
ۛv�Y߆�e�}G��n
���ɷ��!,s��H+ѹ�4��g�(B#�ڠY�O�����#��ٮ������x��J�yC|��;J�K���m�jCj�F��$!�%:K�Oo�,d�_�m���8Wk*�OP�~��z�V���1�ގ���j���e�1}�Ѳ��_nV����%nFJ��C�Xy�0W����V��|�?��K�Is�7$�#�÷
��j�Cu�l���A֎�O �$��5��c���=���������f�r]��p'׎��!�����G��խ��\�� �����a)����g���j�}>����@���jyv��&C@9�_"�;e�Z�;���
�����6(��D���5s	T��&O��f����;��/є����D���lR1���a�!)3$��k��WY�.�El��#:X�gH�r�js�����_��ciMS�^2M&�+6�m$S`��/����k J���f����O�<�6sX�0���X�#�!�	�	[z���^-�26��Dw8v�
!��ͫ[��s{;��J�m%��K���exd j���fq	�dri>k�4[R�c>W"��s�-v��3��i��B�b��[�r���IFOP7W��,����F�4J���������g�)yUjW���_��a���V<H5oܩ:b��W�W?`RFg�b��2Ce�2D9����	\.��xT��-����6�;�u#MR5�ƍ�����hj����}��,�����7�{����Ju��#���]]1lZ���/���dt#���P�F��Ȇ�V�J�x��Jc���<��݀�ͪ��[��
��Df�c���P 9x<�I��<����}�48�Ӝ��s��_z�w =o��r���	����.�����W�<F~na���c�t[��z��.����&,<�F�nU���y�zl�=#F��/e/���)I�� '���#(+�C�|���A��5nP'Y�"<9���XJ���םJ(�c���h��d��" _�k��6d�p^��σ�S\�p����1~.��jٹ#P�~���	������{��7էJ�{�� �4��J��%�ӎC�O�i��8Pb7%s�y��4-ȱu9	�x>����$w/��Ji;{��M�E�̘鼴�us�Q��4z	�H(I����z�a5��"�ޒ�������v�G�S%#�����+���av4Ѱ����i�C ��!D \$�����2D���1��M�]ا�*��f�B�fv��R"� �mQ�w|�5��T�u;��cb/e�Z�����s%C.�U��$�����; :}�c�����x+wq9�w!pH��n�o+[֒r�	t��NP���8�o�u�AN�g=����7��R ���Og�a<����6F3�Z�ɶ@=%�B���z������XY>�E�}w��{��vY-_q^��tv
�d�M[�]�{�R�λ+o!�K�JO8B��S�V���4��$��i�I��,er����7D��a՜�M^_G.�{֪=@<β���/��Y�����	Wx�e��~)b�%����$:���'�.���x���-~m��.+�u{�c�x2Ȁ��#N����*��F�J��,�'yzۧ��$ld|&^͖c�*�x���d�Hfc��aPh�U_~�Xڦ�O�����~�S�p��{�m���wfa-b�J��?���-)���*��?a]���߲c'Y�jH��E���Zy���@�4W�BS�$8�?wO;�X���+j�t�d�n�F��-*��$;� ۼNB2}��eGAMz[��\ϲ��W������;��Ј���uT�i�t5�f�t�\(��������ѭi~텠8J���Z1I�]�}�Q�Āo;�Y�o�_,M#����B�
j2���/�/�U���㟄����ŷ���'璾��J5:!���!��b��j­0pI��uL���3�o�b�����r�Qa��w��A a�1%ղ����H:a�f���˧Pw�>#P��}!�(�p�_gb7�'
a�z�|�ೇ*d��ڏ�r��z`�����(%rMќ���T��Հ#2V?����B.Si���+=9���6<�v?�(�l���݉�ymȷ}�&�zK|������t�`�n��~t�kg!?7Vz_�P&�f��
g�� #�*5���j����~�m���wǹׯ��g��V�����wlN_)�  �Nβj�Q^t&6�1}�-M�9���QaLC�8\��P N�4�{�|w=���>��ȨHUm�5�(l��<�O����=#M����+�P��z�?$@�¿cm��>Ψ�_�9Z�|h�.q��bh�~��|����⥚����rY{.l�k�hPAp�~�<D�k�EG�7��Ε#|�!II%_^��@�c8��*D4�fۦ����t�m��dFq��a�z�k��1�n5��:��5����2�8��;��Q6�%f�u��X��qBJRI�\�e���+o�|�u)/�G��4�`��JZ��?�� ��%�o~;�Xi 1-�&�,#U��(w�I���G+��XNA���\<�)xB�+�.�i��� ���2@�߯d�d��*�����{۠k����i�#t�ò��WO����J���%��e�
���ڂ��~a���\<W���'�ؙ���@��9�v��qc:�N�l����k�ٸ�4�Q���^L�ӾYi��\t���i�Qk�1��%�H}����J��ޢ��j���8�1�>3������I'>��*�,U`�u&c+�<����I'ڠ�4ʢ݅V��T��,ԃ(�Vٺ�i5x�B~`�N����Ӭ��u�M����~�1l��@���ëquz�@O�	ُ��#p1�S��B+�Z%xq0ۜ�s
��I�R��f"�:l�~��� ��X
���)�Y��<�G)d	���|��Y�U���-\�,�n�g6�*LY������i��),��������n�ȇYp�o�љ��(�G��'3�1SSy�^���;c��g@|4y��x�K%�+���-��9O��� �LjgnWø�߇[�F���VB0��jK.@�u��O0��������� U���T��ο���OBQ���7�C�'���ssigsO�&(NǙ�Ф�]Cs�.B�y�_Z	�.��u������Խ��c��m�2�շ�R���J�@h<����t�-Z�|�In9��K�)=����|"�^0���(�K�w90���~H�ʛ���N� /)'/��Ĝ艃`�#u[�.���^�0DY6�t)��\��T�zg����R��	��G����L��\7j����h��YS9Tp��u)?��1K���:�o(��a���P��.<He�����*�ϣ��%����P��SA���|�����K��P+]C��KU d�t^�ꆝ�>EK}�R��_x��V�ҭ=�&��U���+5nT�R�RO��p��w)�����J��h���)��6
םu��,��+ b?%���w�r�?Ř��)�G���@tFA)�-�q�Z=���o~���P�{�f���bU�J�P��D-*a>�O[r�X�:�4�#2��ۃ&(|7�ᶓ�o9��:�S,�w�V:FCs
�\���a�hX��y���D�Э�6J�1�=R8��`w0BK���d��h̡��ms�(�Ŵٜ��XΣ�տ���w�;�Ezk��p|���,������#�|��S2����� |)q�����菺�oӶKJ��QגoLJ�8klq+����1�3�8&E��q!ixn�����sZ��ϫTË_�<ly��? �n�X���`�BF��Y��}(B�|��j�TTuv7ۃl�c��N�� _���HDݤ� �-�T�#��qCy�h���⫺jV���
��ٔ⁩V<�����A�R�~U�]G���T�X3È���O���OC[ޟE�?n���^�GϿ&�������:����0��~F^��/��迷ri�t�v�܂��o�i�ll�e�ȵ2q�#>��yE�#�;<�"����;@>hW�!�Lj4M��p�z��~+G'�`�6�����5��;�� �����O4��t�K�$�]���_g�(����N�k��a��4�kbX��c�O rD��Yx��tI��n
��t
��I8��c�q�:wǊ�f�����H�xY�����O������rn���خ��4����ݎM0�1q�\�vʤU6��o�Ou�[�Q3
"�[�Hu��3��9K��b�A��{��ĭMw'8kH�W0~Ỷ5�5n.4N�ב6���p1e��r�
�&��7���FT2�U�v���U'+��$���%-̮$ՄZ�BӺDI����Y���Tܼ�柲�Z+\҅�&|�{��\��fց�V~�� ���V�C�Q��3$0Mv�^��`�w����_�x1�5����KˮK��[Vf0�a\��=q��0R��2铼��d �lYM�Mb����¢�� �ƣ�/o�^d��K�o"6�.�����ĲQ�zt�њ1�aV�zB�9�����ɘ�}&��=[�FO�O����B$�8���[A@�!+B^Ɛ��l�s��͒@r�9���T�w���rG���q�j�Z��E	���N���eQR [�אr��z#��k���:��{���@ݣ���q�Ճ�3���&� l����NC��^@��ξn��T�m�����5�X��k��ÁxwM8�������������@s������a��u�\���}{`�Ԓ�v�{3����E��M���x��6�*�ujS���C�9E��v�kLj�Z	@��KMHy3A� EEc��X%e�"aa�ˀa��\B_�^�����au-��_�7
d�Fn��v�(��WR��K�	J���`=G�!ʵ�*�r�Ev3���*��g�
�fCwQ]�A��4��-H�+�"U��?����:(D�&��L.��L�x)�I������
�X��]ȇj{�\ۉ��j��8��κԹ�B�Rı@�?��jHbF�^��-����d�þ/�FmSV��L���vv�Eo���:�x�u{�'�:�C_݌�Q&����=H��y]���a|�c3c`����tT��%�x��o��8���,�S�a<�nY���9�kd�n8΄qU5��u<1��r�����H`�Lsys�7�[/�4K�<#�/�»g힤\�����0#�UF���6�@�<�Ge�XW�v����.m,|�a�s"�/
���b���T�M�3���@�>�fb�]8�Ge���r]��d|r��{4��]��I㻡�|�$umH��B�܀�s�r��՛ �c�ڮⲵ=�[H�-Ю�d��&�F�o��:h0E�I�<�x*	��4�Sx��j������Ri4!�b7���졘�0���T��Z��I��\ʦ.:f�3����׆�r�ܺj||z���p�x�r��Z��M�2FC��J��3��o|�T�_�&f�J.v���jv������n�V�YP�_�y�L���� P�0����b�Nj�����t��l���؃MT"�WZ#�d��#WE�֦�e��B������X�ulE��C%�q9����B��������}�h�,Z�o|�A]~f��)��|]�� �Hmd�7���I���|��q&������N~�����RD5?����?�6��TR���>����	\ ��8�8��<��sу��� ʘ��aC~;s�1�)�\��.�_�Z¼�;	mc��{��|&�%>�`�&=�`�I�o��'�L�`+��ΦD���B"�a�/�B����;s_E\k	|�2��:5>LDI����A�Y��H��pM�v(�\K�K�2��Lߺ;���=��D�Y8@�{2�O�6�P-g�c�â4=ju���`KAS� �V�'�֤�b<�x��P��IS�8cyv�Sʝ7@g$r�.aV�{.<��5�P>�{G�Q,6��ݣf��ySuX��?�N�a_U�2����B*���>hu\ݞMwJ:^�8�ڢS�[hE�����9.W@ۘ��H�����}V"�1n�~4ˍyP�N{O��?]}���2������\�l���� pb��X��!�a���*�z��[�Dc^���2��O��G4�v�.�������qU1�v@���[���--�r͹	���T�����Ք�1+��5a���54�f8F�M��O�1�P?��!�[�'̊a�4�5���w�fh���b�V�>l#T�����UD�E��)h^T��3�^��%L6M�(l��^�i��O4	rUz�M���zA�ϵ.T�U�%c�d��6_��g��I*�LWb!��.&��#	m�F1"I�I�	�P(4�{��� ���Q���^�7w���tŎ�T�<�6�֙�݄p�.�jW �J%V���1�
�Km�M�M��WkNCU����uЦr����Wp0S��ۉN�O#�$@/���GUD���<�����e��G*iG�B	+��J̖@Q����=zRhq@���Ct�p}b����ky�ɍ|J�8K�=o`�'"~A;�|��� +������{��1�R�F�x�o�xx�ۖ�lB�&��\����,���SHD�6�掗��V����[��/j�؜U��Dٮ}�˓�s��WO����`e�������>k!�:��5���'.��X�y�����8�OJ5c�b�F�a��DH��M~��Q(/�O�ˇ�/��,�F��g���������4�	���("��!�r����v�2�bi_~��2�@�h
��O8�x_&Z�y@�HL��R�4^��;�``��9�8�_H]���k9T��e2�6*�7�Wq�����KTZ|��G�/&�8�\���7��!H�ho�.��.#E����h|�2	-˸��׀��<��涖Yǡ@P���ɸ�������I@�C�Ɣ([���A{���om�fR��#~�o+�eD��&{�����=z�}P��H�rl��7r���%8��l�VLL�[�'wm)J��اU`��j�q� �qd���'�;�-�(��hݟ3�������n��5	��X��t�:c9�g���gu8[�?w&~l�x�j�E$�,�@;�	��9�ŪGƲ%?4����8�qB�~�\cB2S�����G���=�����_4��ż�$���c� ��1: T��_λ�� ��nslb)$}#ӿV,V���G��]
qؑ���i����R.�솑F�)�!I��i|&�1��f)@OH�h����\�@>V:���NP�C|`
�{�Aּ��"�}-YnC�����D�X�G�}�������	<B�o֚.i��a�������P6	uҽm�깙Ǎ\)��ps4�z�M�iZ|�#��8��3���Bm�觯�_��{��jZ��^Q����R��2j�&G4�����4�{����1�.eRyS�A�5U��]�_���dĹ'[9b��3�"���ׄ��z�*�Gn�DR������%X� ���g^�o�4�4�� >?QJ������I�S�f\�W��&�KS�i�}��v� 6�x�ɛ_"�+턃z#�+��Ai���N��}! ���<���i����%R�ԉ�m�Q�K2n����c/��Ũ+�^y_=L��w�U������cc�'����_O�Q�L�x0���o���4��~(���Kb��7;�=l��� 9g�}�T%���T��q���C�q3b��u _�-�������Qf��pʥ	��gM12w1��ͬ*�ꪓ,�K̄͞��S �+�@ۇ,zS^j�6c-u�g������w����QPs<���rA�E�>�̹	�>H��5=B{n�ʞ� $n���TY? C�cc��c]�9ձ��P1��� "k]�-�V\�e���~:rl�b�E�*�hS��v(rW���+�Y�\θ.����[Go�H�/���ApL����C�s���.Lfd��
�pJA��1��㍔5���y��:˼�-��D���a`A߃�z���yqor��d���*�'�p[�Ԃd%��~���n9��ԕq��z�N��U�\�M5)�'/q���&_
G�e-I�p���#F��G	���)��J8�FrO!�K���nҏ��>K�D�ٻ������ų���j������̀� �n��w��0	��R�6��z��9�5�b<��g2�,��K��.�����؟,�T�9�>vʹ�܏)�]�H�mOz��g ҋ*��{��Inʓ�)�t��6
��T��p�=��R��V���3���K[�������*��F�}H����.3�?���q��{�x�5�t��Gr����ή�a���|"�OF�ļ��qcV�e��h�u<����~��(��j�q#h#6Wť�`s��Z��mv�ܤ:�����j�Kϸ��@d0���aՍ͡�y�7A���ʮ9c_���������#pEMh�ӄ�K�+�PG@!ζ�樱�:���-V:�����,Ysׁ2)+�O�?Qa�߇���jx�p��L��$s%K@+���6�*A.b���^?qy�"�O��b��&՜D�7Ŗ�D���	*�}:O��^�]M!Y�A�=w��z���G����!}��Q�<oi��@�p6)��*d=,րz@B%��bQN/��˞�s���y�}����a����y�Qx��W�5l�|��ѥ��8Rw�ۻa�Djzя�%��t���������<��[��[+IM��]H*"Gͳ�ҽ�5�.����:��;�/�qs�[�ԍ�v��ݸ�	j+��,�V��O�*q��<Z�
��ã3�0���,'��{[O��-��n
�Ӕ5M���Da�Zr����q���#�F5������{�D���$��ds�\Qfڤ��=�м���ժZ����
op~"�Q3��DD<��=]��ߎp1���/���Ӱ�K@u��NW�1p�(�Kx�hTz����� ����.9g�8��~�����gu<0Y�m\��ēu�O{D,_'eߊ�0j�!�f�=ꇌ��lZ��y�d�`��XN�.j�PR��6H0��I�bA�k��^"o��x����I��?<<ʐ�d�N �Z�Q$ -H����83����5
@r1������q��l����4����-�����ƻ�,�$����`��"�,X��D8ZO����~��i���)��=��%�r��$x7��s^%zЛ,C�1R�a\�}�g��lc��Ra�8������b��<���(x���
W�r��18���(�U翯�Vw��-�G�����L|�2Ze�r�c��8s��P=��՛|��E�:����ޅ�叽�Vye��^Koij=������Ǟ�H2x�!�|j��{���1dQ�8�~�|O��q���ǃ��N֛PEi�F1��'�[q�2�BR�5�	'5q�P��d�D���p��QK�_�>�_��.Y��P�M�)��3>�����T��꜡m���B�+�p�خHn7��R���֮��W�gг��1ꄸ1[S�e�Q*�9Q��'��$A��+´'D�D�:Xa�e���D�6z����/�
�2��:�@n��P�D�&�Gg3b�����]�b,Ĝ�pծ*$���䛸��7�FmE$�P,�c8�¯����Y �CXZMQ�`%�mJ�LœWT��>�O�$���"��#�iGm�ˮ�����^����iu�����U��xT��#$���L]kuɠC.mYQ�jRz�w������<����o��m�Hi�"��{���\���1䰺4q�]��흄�5(@�����4�Z��+��ׁ�aB�U�)��>x��պ|�+R�뷯xR݊�CG�`���{�Wc_	�0�+Vư���q����ka�э������
��9W:���'��9�LS+e�P�����L�rqŐZ�IKy��|�	�1����I�+���c~�tv��z�:c*s�ޭn�0$Rw�i��v+��%O;�^q�ݎ��PG{�2KIC1"p�E�*9#����}*�U��i�H4�}_��[C`m�j3����q�$�Ǌg�a�E�=,"�j���o�na���|��be���!Ю��ItG�v4�g�2����)�4�O�F�`��E�E1,��X��ß��Z�_ȁ��Z�Mf��w���>��aa�����$�*@l �G&�ؒ���^;n� ��!??���h`AqSv�tnxwm	����s`3f�'s/��R|��H��?\�Q��\�;~eC�-z��+am���y�_@��dY�h R�թ&t��Ϧ��/3���.�Eq��Q��Z`��k�:�H"�+�7IsMjO��qݼ���?�Q?h3ֽ��;���$;�.���Iׇ��ؑ�dADm�����g��㕓�����'
;���1rǥ�A�����< �����[��k�H౶1,hh%�+*���vJ�����Q���xhb�2BƯ��N�y����1�4�4mE�Tw�H�ΡF1�fv�����	
2����H���1��Y8o���5�=�ɔ�	� ���>�����\fE�X�;e����N���+%Z9鲪�i\��j�#����	�	���le�WҮ�mtb�g+}��7z9�v�QQe�uS۔!�!^�+�,�J1 ��yǾ����°��l��S��mE,�'�{)Z��"غ4m������h��l���6'W+�&��ˇ���z��?���j`_9Eh�W�Pȝ��0 ��-�ݽ���;d7�")R�#2*r��ބ6آ����J��u:�!��zq�%Zt�-�s��`�ޔ���yRVC��4�A���r��"�������e8/X�^K|G��:7���ُ��6{(6k�o	"��e`���i_q?n@kIӎ?>���Fų|�H)�����L��O���Yo��|��6/w��؃)g�'�D����-�	R�Ũ�t�>�j+��,�ؿˊ�_�	5�I�m5���ar�qD�����M���$�a�(�U�{I޻N���&�f߶A�(3�9���g�N������{�$��c�wl���j٧���v'�ny�{M�J��]"��:�{L�lϺ�7~H�;y��������b,EX"d�[E�?���ѕR�C�ţ�uDXx�,Zt��V��`��ڲڬܞ�)���%W��Q�}k(G�V�:�2�4�6�����nk_QYԋ�<_��$&�=3��}��3�2�������ä�~��F�
�@�@
3��6)=���X-+�g��)�����>��G{�ƒ%���+����>D���N�P� N�~��F	y9-=R_�Ɔ��5��:~�4����9E&�?>�W;t�",�s `\�Z�6XXu�&��>c���&�O�21]���<�f=N�:}V>��'��Gpn�}O����e���N���<�K:OJ��4��##�CT�!n- Qh���ɍc
!6�XS��B��s�n���HQ�7$o�4��ۋdP������u[��2�h���XV�w�  ��7���r"�9Q��JӮ{EIQ����А;-�q�1��m�A��!$F����K]׌7or�F_�@$��|������� �o�-Xވ�:`��ވ��	3�J�QNngc���BzV9���b*aBB��L��L>^������Ӂ�ۋ���S0�b��+����,�~Ї@7�gs�)^�[/��E�ԏV
*ZBp����)0`���l�:z�T�3�~�x��*�lu��>l� 1�S@��UK_�mn\��y�m�{(����4QޮJ��P8����!b��Z�����IC��6�bZqg�к�Gl��@#}��肜i,8i�A���)Xv�Zz��V8�,VT�ڕ�g~âj����Jș��g�G��`=+���qe~��"8� (1�:��%�-��h��&�W��L���9�4w���5r��+v�<3��=L�<X���Y�eӐ�oF�5�� q�$J�*���s�#`�l��Jd@C��	A)��<�p��K���{ -��'hF�i���H�rf��F��N0Ԯ��ges��ye�ULV���~�V����?�����To�:��>>�G��ڎ�d�}���iw���O��U�'!ѷ�����:�CmsC���{�-z3������&r�q�G|�<Gf����ѹS��n�IV�\����)�����~�5b��u�t HH�R_}R�j�~ّC���~4}<܃b�� p�q��9o=�cT���ơ�� #��:,C`�:���>���+�i;=`�3���}��p�e���Arm��Y�{T�ؿplz�T�T]?��Ȼ7s��-[V��ǴvǛ�]�?[|4O�_��ȟ�U`V젿B�9��M�[X��`���Щ(.	����d���@�Lm�d��[}���z�t��:�&[��?"�ʙ�M�r�s���Y��oZ�0o?=�j�5��7��~t���b��k��%�2ꕎ�4~�y�X��b�i���36l_���3���a���%G�sݫ�z]%t����ăH�.���P�~>��E>� ���~LŹ�:a�c]�g=LȄr&�;����t�(�f����;a\��ך��_Rc��3H����1nȬ1~�b_��n�x��oԢ+�欈uwJ�)b��0Sꍜ�����>�'yq��[�Xl��KU��)���xZ\[�m�Ɉ�D�!jw'��e�J��ʗ����~T���bB b��%	eC�Qm���B�]�r9�S�G.����̯Q�����r�~L�硩҅A�����zĆ���H|�/MӲ�����:CS雎ር+�p��{t��U�'l�2��	�:!� �zB��Oջm{v��c4��Foٿ)W$�i�W���#��x3� $ZB+Y�~�}��k��KZ3����ف��6���� ty��v�Em�^]�k���'�}f��&$aE ��-����M�'�9��3	}PΓ�5�T^�S�	���a��]7�F�+W�t�8�4R�GOȚBR�sF1<H/e��z�r�:��*���wC)1S���$�뻼?��<����týA3u"�T�w��x�<��h_�ML+�?v�"-������Au�yz|1��Ew�>�u�f�S��U�s2d9s<i�Ζ[����o17���j~V�`���r��wò�҅l��kZ=.|Wq8l�ͣ�)�b]qcB�a��m����KW�V�=f�YϮ`)ʱ��雿���O�Vy��r@��Jm1�����@X��eB3AG͕��#����tk��jO>!�#	i����-�I�6���G�5a�%Y�=,V݉�)�`��v7[�����J�Q�/�?��m�#����1?Ukt��!fK�T�+�I��a�~���}"���n�NM��j��;c������)c��O�Ƀym�G	5s)5JA۪�@#��Dr2	t���Y��	E���n��#h�N/��Ն�J�lڐ��i�ꦜ�C�]�����Ӫ��ʈ	E��6�����b�9�\��y�M����z�-u���H+��"������6	���|���`�)��z�����!
 �]�9v[)"�XR$��rj�a�7�C��g`]�,if����1�M\�֬�F[q�l��� �%!�)}ώK �I�a���ψ��-P�u����]l�qt���8!T�r�w=����Y�o�Z%��$X�n7�����Ս&����0�d?���$o����J�e���+�PC��!�����n�5�f��// �Ň�P���[�������'��$�7?�SS�Rs���lݍvWˡ	�*솫.����0�'���~�]Ǳ�	B�*��O�.��_�bT��<S��H/'#j.�XR����LÃkMO<{B���!��K?�pm���P�b��U(��UA#�!lj)ʗ亶�_�Ak�ҫ/)�sG�� x����<g{���0R-0�=��0��$���y��h3=�q9��Ce�4������3g�����R(�G�^�P���DXX(���ns!�#gS��Q�4!Q�FL��トd#4��j���0u#�F��g��x��/�7(S�e�Ϧ��,�����@�v���Xm��8��E��H~�P�ݤC�1�6Y��|׬��3���$�H�$!J;."�O��W^�3�"F���>U`������!��`���"��4�i��S�ؒ��2_�)p�h����Ne��ȅ�9���'Q�����g��N.� �8�;�7�#ں� &�������Gt�b0��.͍_��`��P�$��k�`y0��*xv������:K%���z�?	>Ц�=�©���љ�2>�'s�W�@̪�r& 5����a={�#�0�U���h뵬�+�U��l39%p`:F�n!�|��Xs��x���`%���H�\��Q.	%:Yo�ʘ3���:]��&9��7x5�Ş7T2hn]}�Rä �z��j$�ßTPNK�F�t�&�9�{��{G5Zmq��Py��%��{�I���y��ޣ��$��s@�P�zܥ8��S=�a��Sez�l�8��T\�~o�ޠ�t�m1մ����K�N�
���B`�Sq��[�h;����D k�0��a4��UE$��A��&ۙ�����j@���¬�����K��j��eq��|�Aћ�&wŜ�68��'��LJ�|I�FU�%Y�?z=s��5�Tx�>��,ΑR���|���v�o��m�}�����p�[�qE�z~�3�n���!O�q~�	4'A�DiT��W��A9��\�A�a>)�i$��|'ˍ�za��쩥�ҪE��y��#Y^��-7�R"Ҡ�h��:��3��Q4�aE~�&j	���Y�<������J��??���$\)*jK�6櫝E�+��G���k�Hq[�(a'�d{�B����@�{Kx���]!II5����!&��c�Җ�+��ǒxIc�}���١�B�D�hת�L�i�%]_����k/��=��u�3htG�$VFD�Kxq�3l���(7�ֺ�e�E�-��*�i���q���(VO;h�S�ɝ^�F.��X� jOwgY�pS�:�<��i�rcT=��Q1J�9��Rw�	��^�x+g&����
�CV�_����o��Γ���j��P�F?���)�)(ʱ�| �n�Y #,�]+&G����؎�:�=�n�*�(����`�JE<�)�(�.LV>����j;ltyS���#�-_����3�'��c�~�j�(�E���7B��0�W�T
�Y���;#��G���o��T�{Z0*�xe2�5e>���6��F�1�,�_Q�P;j ��$SH}=��O� ��ȕ>6dqb���0��y�~e*1�f/�-���L2d����$b��A:	��%
�r62��l�I!���4�R�����s��{�( ��;��%~���N�i�=��3�(����`L}�Q�%.��)���$����UuEy�y�2�O��m��=��=B�0�b
�$QKz�.���N�
��,v䣠��������-����A�7��֌4D$��`���\�=
�BۗN�q�4�OM�od��1*�����u��y�b�:��=��cw��Ƣ�!�Iᣯ�d��n���Url�Y]�C���t�VwLo�;���zT2&♗��VO��sn�X䖮`]�o0:H�|>9?����]`̶:l�$<��\�-�,��#�Cq����_��!���`@.<���
2z��]��6ױY4(>p� �9��I��J3����x�*����b�������%=��.�#�(�5�#Ȟ#A��1�%���F�I��o���wk���]L����L� bG$���Z r�����pE5������sK
C}ɪg"���'�@�'p�����DܟA�4!������z�.����Z���m(�t�i��,gF$��������m܉+����I]�|��|�I���N��ǋ��\���F��Z���E������n���dE� �H��و�8P!�V��s�/�R�O�BC��A���*���>Z3��?��ٕW�4Oٔ�� Kg���%����i���o஗���x�嬯�Zx}�u=�y�W=!�mc�p4��)����g��q�i��۷ �,�}mJl'ⶏ�C_9��bE���T's�<�o�ƈ��~�d�6a����ʿ��07~R�5h]��+=�>�یP������Z�pd1��"�.���U%�;\�&q�QfH����-��{�	k����H}��0�	�'���,Z{e97��Y����U�y3<�/��/�D�-v�O)�tZ �m�Npz~=^ʺ��:n뇈5↨�|c��.I��|��C��*��Tv<Z��J��/�o��� =�JD0I$,'tlpj�l������=��?W����:l�ԉD��d�\��~��OzFa�͢%��n[w�k�\⟞�(c���ұ��Gu�-�4���f��t�x��6���g�T�#�R�?H�����J	0�a%B>٫g evp�У��YO�_��3�����K��$q�Q�;����z�g�t~��B M���_K�T�de
�+ߵ���@X�0���۰++{��M�\�-�ʅ<-�FV�po|�~�˿�)��7T��ֆ�����g	c�#*@�|Zߍ�U�h3�3YK�WlPy��n��R#�A�dm��#�Lh;A<��}Yf���}�,��}�r>�Mg�Q�!��^rֱw�����!�S5<W����>o���&�ִ�(�g°������G���߫C��e�$�L�j�[��W8Цޘ˓A�K��E'l���O��+O���ܳ=�j���j/�?���Ʀ�[�������גh���Gl�ȉ��R���d_
j�-�8�"��I�#<�ER֛�Q���s�l�E9!2��8����(��Y��:�9�5ZN��B*�,�Ļ���7���	{�� ߆)Y�#��x��8?�Ӏ+���cپ_�*�,Z>�JoECd��rֲqm���'HW�?]/Bg�9�����(j�w�����ö㤿T��U9i���R��!��ޡ�
�^�;����Kw��J�71b}����I�SA4�C��S�!���o-q�O#�Ι٢�x<	��7�,2��,�TＵ�1V�]�\�ý��W���R1��*1�8����� ��b1'I拙&�G�.��V�ӚLQ?���F؊ԶS���W���?���B����L�c�}N�-=���zk���-� J���%�a������@-��`�o)Rg���1Ώ ��|��.ĤUҽu���%l��F� ]���2=�rhl�vI�V��\�nʅy=�|�ȫ��\~�>;a���E���[Ȃ
D�aF����v͊�e��E�q3k��=�DIc�֣3��0RO��˂� i�4X�E����M#2����+#;X�TN�7�OF�̃�mm�(�h��i����H�c�ݡ��W��s��Fk�m�0=���KZ^�ENx�����WЂMQȃ����B�ː��_���0uW�����?���!I�[.v"�sV��1� 7�3$N&��"tn������k5�Eq���X����M�p�kܙ
�-�%,B4Ccw�U�G�;Uh����)-g�*|.W;	⚔V����j�+僡�j��(��l�fT�u+��hą��Y�{�]�]��A�YK٩P��T����x���)�1�?B�rg�M(�ŗKR�X��#�Zɐ�����^�7��h���+ۡ9VM�=��\�19����6����� ɻ��߸a��G��n��v�C���C���������V��[ғ�|b�.�时�tB8��PQ�<-��Xd�h�N�ZIO�j8!7�^v��x���OtQ
4,����S��G��F|?�u��.em1g�<<�E���*X#��.y�X�s�-�x�����l5�(xbQdV�)4�Ԥ�Je\��H��v�W���/�ءC@Fk��*
��m�9V�.�U h�($s����ƿ��7�'�X��������g�$�E�&/d�љ�N2�GOT� Ú+�K��m�Eb�ֹ�p����^���S���q8X�q��75�ܐ���~V��Q�lH�����M�ҕ����QzlZ���7�w9�|\86�����r"TM�Gw��~4u�-W�x'-�w)Q��
=��\#�A�x�iɝ�Pˈ��PKD��3���~}���1p��#q�,�칼aZ(-�co�_�P�Po��g�z2y�c5����m��"��Z%m�d4��ȝ���=�vH�X'ra1J��a�b��2��o���9�<b�����̥�mgWdݗ^�~�e����z��Wi±��?�� )���Z0ſU�~d���r7}K�}gRci��0�8H��V2��B�-�z��3xfX����Ww��ob��Xf�z�n�n9Z��X,�,��K^O�~G6���`�ŰSrn���j✟�1t��	�uƯ�1!�#�R
;5�b-�����:t��
H�`6��A�9�gn�Mi�P1��%��<�����R�(e��*�ok�(�zfD8-�!� ݜ�E��v��{\���ӭ�0����r���rd�)��?B3��T���Oa���O�-��J�H�a,ۓ�Q����_є�d�������&�0V�������Ot��-�W�_�Ƚk��z����)t�@{Z�	YdC��i��L��î��p.n1'��_�2����h�lK��,H$5��e�>����o�z)���E�0��(���:-8�Q
w�+L=��F�Cb����6}t���7"�t��'@լ'v�]
��:[�^�P����^>H8�nb�4\��~�4QP�L.��H�򄤱�~WK��:�=9�*.B�6`*3�[b��s��]l�k-|`��Sy6J�$�;�	��\$��^{�Y	��X��鉻��k���J̠����0��r���	�Ľ}#��Xf�9� O$�`)�Հ7=2��6��06k$�#���q^NW��b���N˯�IdB�z�M[`�*��Wn�w�w)5�Ɠ�&�F�	w[�F=�~�u�z��p2� �����7+�-���#k����Uys�ʺ{�x&�:���:��"�X��y�g�l^���D��_jt�2�_%N��6��{��ݰH42?Ÿ=����X؍�'zq����iX^k��m�)K21 �W��L��Z��:[3�3�]� =}�e�JK[ ��վT��&5*��m��S�:��c�����N��{��ǯ�)�w���G���<C8��>�~qi���������� v�ҝP����b�X|<oOc�h`Z�e%!#w�d���,j6t+���&쩠���A2nke����6�}�q�M�O7�t_�`�ez��-i�
���m8�u�ٴ����~��/��\����'q�q0��4�����a��);��FdiV,Cs��*��y�+���"L�(풗1����� �g���,o�^b�[PRh�,+��W�642H'��AṤH��fH�ገ"]  Oa��N���]e9����*4��U��v<'��'���A��H�Ɠ_.r�a	���;�Ex��R@��iH�A��f�	ܨv�v�X�T���j�#�E]#�P�)��!���0̫�S򫜮�&�����5X�5��%Xc�[ʬQ2�������2�c5RL?�<;�S˦�UwF�Hq)���8M�\���7�g�����Z.RYMmںJyN�5��*6��9[�0x{wC�z-Ɛ�����Bz�Mh컙	2(�-�?6��{���ct?��ԋ��d�ֳ��4�� �Un>�ƌ��SY��S��i,�/+��}��6�AwFI�^�`��
Q �&E�_ʆ#Z��vw�q� o^�BC��"J�g\�-\N(ɢ����(�?��~����$I��
�?�'�5�K�P���^��p�ӹz���8��_��G�7	/|�A���	�{�g{��`]�c���s=ݘ4 ���}f5�Z(CҐ(4��j�{ *��jʗ��h�� b�t―e��`�j�#��Ph���M6߾�_g�����v�e���1���!.m��KIp��YX���z�����5�@����G!p��3񟵐&���m,�R�̥�%��6½K���y#��)ލ&l�9|=�5pdGm��?3��}����!�s��~/b:��>���h��im�}�#�$Oߩ/~T����+���i��:�7Ԭ���3aL�r�hb�+��^z�e��F�&t�3����Ҳvv<cw!�P1;��%�qs����v(d�\���]*�RDԋ<1�!S��!'w��d�\�V����v�);�H���x3�`�jd2��P\,���T�ۯ���#kZMy��`�=9�t��z�ڬ��ո1��c�S����X�"��J=ni�
i؇o�ʿc@1��Ys�m�J]�8f��paE4s0����,Tt-�
"�%\�L'%��be¿|���w�UD����U����*2�\�:�ݴl���A��.��o5!�6	,Z&�>�3#\(��dK������F��jQ}�]>��V�-��:�Oy�KOO-��H�Zb+��N�_�Jf�]�gU��Az��ȧ��s���3/��`a�R��-�~���A��V��ږ���
OzC�i�C����}�gLブ�0�{�`i��\ǥߪ� �t��,dw�gH2�bR�\�\ʷ�3N�"Ⳁ��4�R��-R�o�ɒ;�,�/��"���l|\{R6���������)�oP٣X�t�c��h����0����=6��Y����P�ݤ5����rY-V'%��	�S0����@��_x�f���2��&�ZI��b�{J���r�z�cĐ768Ύ�O2��W0�;������lE��ٿL�������-t����dl�د�]�d��a�Fx��\�t����Qeqf�g��,I=�����x�[h��8��J�[#U�?��iJ��4V+�td�y�'��-t_�ir��,8v�(?Q�o�t���a��@#�e���izA��������~��Va%���0�5b��j�Qݾ���i�N"����	�)�.�?��ezo��� �Of���S���b�អ�A���"�.���O>#Q�Zv]Șh?�=;8m���,�.X�~�Os��U{\T�,٨�~�n0Tcɕa� q��Hr�ۄ��\���u�v8���M�����f��	�7ߌ�#�[2(������9�ւ�	"�%�iP~$"��j�(�X%8�������������c��被V��+�nL��ʏ�=X��`�pC�}��y��]���3�!�
>�]�H^`�A{c#k�ʊ�������r�ݹAk��S�}4^Jaa+��EK����%W��L�Y�+����M�<�)�]��%�2�ʾ��ǗA��`A�?���SH������HN�Ã�܌Ao���6*�@���[{ �E�'���<.�w�,�f�2&��z)�^�ĝm�t|KX��I
O���=�;�7�3�_Íٛ����Q��׻�?+$ԩ�� �=��}���<��Ncࡒ��"J��̖^[�����n��L���C�㱥���_-�ڶ%r��HE����<�x�U:�Os��E��=�������led��8|�B���v���q/�j�;9R��m㓜%)��eq�ap_St��;�\�Ml>��>}ѭ�qz��pV���	�~~��<4�ן ��?�҃p̓���|~�|[��kf��P�p�-��ζE۾%�n��΀��4����5W'dY��^�gB��ą�&<o�Y/�d?d��m 0x��ZwEj�;����|aL�����Jȋ7�O+U(l8U&��6x����=ӽh�]OZ���=������V���D��o��R�e��YYډQo��`Q�Dѯn/WK֧�ಊ�8ÏA��
5��"�d2���K �(u��#]�v�G�*�~�X����1o�ȸ���֗ ٫	�s�8�|L�D��:�9tu�=�=�����6�M�g �N�*���xq�������&�����ˑ���־w-��g�H[���mm���*��� ����&D���U�k0)b��c�ԓ�� ��8�Ǌ�&!��eqf\b����t�F����K)�06�'�E�|%�L&�i�0�D�K��
��1"�.�r��U?e8��r&���|F°��Ru_���>\�QЦ�4��S����δe�?:�}�Q�a�M3z843u,O��}���Qu����QQQ�^|�f땄�Y�C�x0�Z��A�{���4���X�N d}��7��`/�S�P��)�F4ڛ�,����>�L�E��q|��&��<��[* ���
��~����h�[��IĭHHJk�ũq��ez�m�����i|@Ĵ�X��o����
L�Z�f���$���U�p�4�7�+�:�kϛ_�k)�L�t1�M7�f�8��ʅO����	�L�E".n.<+EJ�e�ڵ���9����pA�طɨ�+����K�3�\��������ㅞ`�ޗ >�r0H?�]���z�
���e��cg��R��9\�Ef�3厽Tg-���h��y�۝���.)�������x-D���kD�X%���s�.�TH�>f�ߝA�)N����\�Υ�Sa�4��/�A𺅈K�З�g����B���z�����c���_ޣc��_l1��!�Y�Očh�FjT%< V�5�lj�,���y����ɷb�x�D���qK�>-�����u��J����<f���{{��A)�{��]c��!�QR���R�	%���.B��5v��Z���<\�4��_c"���[,�:�ۢ��,���u��njT6	��x}y(=i}���3^]���m�=��S@��>�"�I����G�j3���0�ۙ�B0�-����F`�k�b|���M��e��L"�^/{�3�"�Y�����e�r�tNc@-�Ty�� f�8$bъ0}����άl	<��9S�h��EprbF����y��ML7$�q�S�a�5n)3��������K������d���
�r�u<@�
x$s{�f&3�yqٔ���9Z���o�*�D��V��>2�e���H�s�4�� ��[Vѭ}�	��{p&��f����O}�D%��#�&����uV}�RW��fI��d[�8 ��Y�P�2xA���&���]�kB�7����'�q���u��P��x�<q�M�1N�^s�?�*{�r����uv\��߻K����l��~�9P�d�?-�i������F�� ����t���'?>o�a�{nM*iQk�9�2,+��tx�]9J�f;^Ӳ� M��lbۜ�r�y����ф������5L*扯M�V&�?vuo�L��%)y��������es�a��~(%���T'9w�����`2��M��u��*Όb6y���m@�O�H1�j~�3���i�8;
�ۆj�d�v�N�/��
�j�a��%T�,'z�S��4,�m?E����ݠv��$���P��ȅ�!]�l�V������Z!cfׇ��-w
��h���wOYJ0�4�S�_��H@��S3=��
Jҕ��E�b��f�z!�o~?Cj�����Tҝ
ij�7�0fε��/f/ﾊ%�kѕƤ)#7�:&	�?��Cr����ź��1b��^un��7�($�S�Bul�L��fJ$Ǯ�@4�X�LS�.���v�K�U�G�x��I��orkߦt���Y8��=�����fN�V�\Rd&&T�t�BWen�T#�S��o;`h���=	�(�4��K	T�6r^�0��Z�W����Qrr �E�l�OR����~�A�+�\-��~���ajLg��S��,$$PlU�&�� ���	�<�s;x�TZ϶ٸ�tΌn)^wҮ��X&�tl�~��R�����$�oz��"�\�Et��ކچΈ.���/|�̍����w��f��؈Q��kp�kS��<r)L����6�nM˝����<��"5���vG�"��m{��h�;�?L��4(k��Cخ}t��C�b8r��)9E��D�j
��\�&�me��Z���n%v�G�F�=���jn/�¥l�"��Աs	p� /$w{a�Ӝ��}a͵���9���a���;y���Z HOQ����9�;Uf6�c�+�ދ��^���y���Do�6IW�.��Z��3���^���7������0�pk#�(��F��W>#L�8��{-��@"wڙ�PJ�
99ZW�g��GT'��%k��k�>@R�~�P�F{aI������/{~��v9Zz�H�3pr�g�`�u&;�h@}�H��Q/��a�yq���f�l���-7a_%jK�x��PU�5�Bu��8q���̧��Gݨ-0;��[�um!�Kf���3����:�*lq����:�U��3���Z���i���*b��0��Yf|$�o5����w;ם)TL](q�\������`@��4N��|Lg�]f�?C�mv��VlN�}�]&��D'D� **�Y-2�#��v^�Tir�PEMݽ(EEbDC�σHP=Op�2�L��o���� ��'�R5l�3R<;_�L �j%SQ|���!֋n�l��ߞltL�x�����ވ��f�B{�+-�wZFԫ�2�x����#��ƶS���$�#����}=�n���u�J��>�V�j{���w/~�y�Z��x�(�I�)��a�6��K=E2�NM���ٕik	;7�	�q�b���Qq���^َ�_� F�v҅�#]T]� s���)y<�*ײ�$�B"ƽ$���[��4�$|]�+R��}r��Q_�j�+H.�l��iւ�z��n*��a�g�@�S4U �t-)k�z��ɕ�1�x_\bL��L3Z�;���"�ב�X�֞|�+�ؐ�ϯ������z߾��lox�?,_T2���9=��E5���`�Ѽ(7����N�f��]��K�SD7������>R���r��}��Kvh��m�~SՀ6�N�;�������AW�kҍ����=h�AJ�,p�?�b�`�\��-��"��;gN~x���+��ǎ}|-F� �l�q1�,�?H`�\%�����@���Zd��V2�!�-��`�j�&
��T�j�����W%���BG��.��7?�1�H�蘆Y뒎U/ /ܤ�����|�A�t1f��	�����]�Ū@�aj0	�T{!�m�@�v�#�����O�Ԑ�w���n�Ub?$t���d�ps&_�{͚�.�K�� ��2*��7��s��TOxJ�+�c	���(K���Ur��Z�����ш�>b� ��������.W��myp<Ay}�Dsb�[�y<\aE�7a�S&x��_S\p��ы'�v����_c7O�"���.�B����o�jzJ
�t���X<	ۺx�W�h��4�^z|���-��xG�����$�)��Z�;[f����T�a�PL�\���H(<����P3I*���p�GZץV֟ǉ34&� q,Pt�D�s�z�UECAS�Cwchy��O����:g6zM�"?��g�r}��|�M���i���a��%IP�t7.H]��-�dˆ�r��t�v�kv9�����H�8���L����,%Tk�񼵳L&��k��P�k�*��3�^u���?�H)e����m�i�[�<Q�,���&����p�z�PM$���"2�c��l�ޠ�l<�u"z9�0��&#H`
޿wV����|��'�\��\z��k�D�;����>!�E$̀/����d!�o�DH��v�n����{�П��<�!� �%�Pʐ�H����TXÏ�s��w�!�0gvX�0{�#:�{F���q�8^*�e��"yF�%�UV ����x[�M��S�s�0�yP���4!���Zo��I�ǳ�w��w�F�`!�o��~�z��uIS��f�^�+nu�
ݰi��*��������c�o��K-,�[���鈍J�9�2�%/^+w)d��G�
S>?�	+�`�FX�:���CL�DCɲÚ#�pJ-G�*l؞]����RD���
E��N`�K���i�ut0����O��'�e7���j��	>}-��6iL�6a<�s�f����E�h�����B4�=��=E�����6����iq��;}�:v���A��X6k��q�m�:���M�_��aKʒ���kU��\�r�`��^�d�x^���7H���4�;�F�p �<7Es�n�� iU��m�iKl��7�$���o������sfa��p�q��3d�p[!`H�
��A�f�j)�c�`��領,ә���K�X9���t��8��A%��h}�L�3%޼�0K��p�G��r����;>��Qx"mH�k<)�"��3��:j(��ݧ�VƄ@:fy���q�JAYQ�fXm���^��<'hõ��\v�J�
�q��˝|=����"�chS�퀚\�Mw������x���Շ\�����)hD�s���.�M��4��AkKO�-��2�)j��߭�t�8G�)��XS���x��c�2��{D��@��ǰ��D�>)!C�cU]�2*p����7��T?�u�6	��ޟa�`�6�9V�5Z�h׬�h!���B4��ќLS���q�zȺvd#�/�d��Q�Y�%�$��٤�fZj��X��!Li�|���ݩ}�T�R{�ڤ������h=�w����Y�F��u{?q��~a#o ��L�A>zE���) �n�/��c��6�z�$fm��%w�o2�����.y���1ۙ����S�l`��rϗ��	Q���va��6F�N��H����3�*d	+�/"�.a��%���.C<b��l��#B-}��j���"�"v1ײ���!m<1<���P�����6�L#%I�AD.s_�ab�*�qrjY!��]v�T�7'�vϱn�*�/��B��=U2��*�K%&�8�hl���;vԾ&�A�Gs���a�O�|�����G��Y��V�F?R)�J��j�L8aS!_s&i)8p���˰s���_˙s���jMWw�nK��b��Y����03��A���R�p,�pO<X�+6��.yODk��r�����颙VZKjot]�m�}����s:�W��,�)�]sp�Kr>��譽5�ˌVN�~oH�[�� �w���z�k�O���`w�,�}O�����b��y�f�W-Lѱ]�Aґ�Y�q<׆�H�6��>F+!S؞��l.�kI(��!��}G�lq���iu�d�d���u_<�@ꮇ�24���<QUF��������>b06�.C�65�<[����ʳ��p�S���C�5
��}�W6`������ڀտ��4��(��e����x���=-XFnKV�C]a͒���ڦ��*��������#9��?~|��`��������|v���P+�ϕ`�g�ݼ�%R>�+h0\3��I2 ,�q��� ]?�+��j��Q��M`
|��M{X�3������`���fӤɚ�]N�40��,1�{Q�6��z����Y���:;|8:5�c�e^�^�ۄ`I��.2ŭ�]��%l�սȘ��Qۻ�ϰp�u:x�WW��,Cإ�Xb��BYr��R�+.@�k�U�v�򝭶KC�g�[��R���J�ӗ��m��;�������j+ҤE�\}���.S�{z�c�Z��T+XWr:y|U���������F�8c���ek�&/�e����Ce��W��$hj�*��=�F6̯��V�N@��k�}r�­P�G	���	��d��Y��3(�K�_U�T�pR��)���a���X��J�o`/�<��Z`�uM�!R.�����U��٪>B�I���.��$_0�� P� =�V�`Jeh�W�'��XRPg%| #%�-�8nt]����,����������cw~Ƥ\�:"� jAǈpQ+�Ȇ��@�3�i�K��~z
�� Oj9���6�І:36�,�Kf9=삛����ٜ�4&I��-P����@��]�AcW�ڐ0|���xu`w���8dk�k�*�$l�g����N�.����(ܰt��ަ����)����i#�f�x�:��7.
we��k��v���\�)��k��5�S�<W�`� Z���ɓ@ O	�U������CZ��| ?�!���u���.C�G(������-y0���Gh�iE_��;j���`!�N�&f��[W��m�}��B�3I4'��)�ɗ�~��ӗ%?ċ�e�i<#`,l���o�c1��8��6���O���?�FS�R��T��:�<�&�rDu��[�jvu�7�=��12���9��M�')d13��#��O��lɊ�/E/�5�P_��S�(�����ہ��j�,���G��K�6K�Z&|9oOcT'PL�e���_��u.٦�RW�nҳFy��1��>�A����*��F�+���բR�i��'�%|#hmgrC�v�I�j�K�Tf����dS����"�
�P��ҫU��b���QhtE�k��
uu^�g���ԧ?�2�([7|GV�9�g=�>�b򵟗�dEc�Aۓ�w{mM\͏�4�H��BY���MxW޵#aY��_�H���ح�-:�=��W/�NT���*�PD���}'B��/���en��T�@��?^RLo����s~5B0���R�p@�͌���*�j�7�AH4t�{�mY�(�g��|��ˠ1x3����1֟+��;z|&w���$��'i���JBx�/��m�[3l����������d�r�2���#�+��B2���V�������D���"V�PZ����K#?{��[��U���vܬK�_�~�Zb�J(o9{_%�M�d=�Cu������I��T�?�@��j#9��%��i�p�o���:�ɉ��y!��F@uj$�f�ٴÆQ[ nMi�`}���-��I���>�k �S(=�f��.%	}K��u�W� ��F=� 2���h��G�����9,���}DT�}|�\z�\����>�r6���h1�<�Yb���Տ	7�;�m1w{I�C�hl�
ٳS�Z��/-��5�ȘFe���.7HY�����eeH�'!��%LF\�P^1�����gA&�fZ�1a��h�F�a)�C^:'�����7\z���<qn�ՊB~P�k ���[��s=#V������0mZS�z[t�^��_0�.-������J�J�*v��(���'��U;����q��� w�����y��z��s�ۚ_�&e�:5z�±iȋ'y�IXxDP��?�� ���ƣ%�__���H�A�@�����N�!`5������I�D�o1v�P9O�T�x����\TuNp���wo�P�T$���-Ĕq������pSz0���m��&�=Q����Q����r�� /4x�K�؍7 ���]�a��ċ\��L�qs�#D��JS�0!�6.x�[�A2@�ɶQ7�>�-�F��0ڣ���tR�|�����O���r�Չ���6u޳V�D&��{�A�0L�&��������|�]��D3���B	>[R%��{�N�H�K��V��WTk����O	��bi�nP��/�ͪ�{_����c�i_F
�Q>\���_��}�^���A�B�(�1�Z���sc���{���Q�oY�P^Z�h��2"��>�.��\g���P�2$nRWO�SK:ݹ"�ֵ��!e�b�FXyT�j�V1����.�d�o��֎1�?&V������afq�n��9�Z��*��uK�H�7�#>�P��~�*��Y�	�_���l���ݙ�P�o2�~k���&����so�xy@���H�B��0��S��}�;�ݿ4��U��rv{��9�#�S��x9r��9
RY���y����M�8D&{aD�i1{ʟ�wf��� .RY�C�}QnTHAsN�"K�0%T�
�����6}�)ɯɓ��+K�����~/!��p���Yz�[I�H:�`� �����)	"�Y�(�J�⊎1v]^r���@�^��L��|��)�d����SO#�QC�������{�r>��>+��U^��G��<��`��T$a�Ue�u��Mmq�UK,��(j���TZ'������݈ю�Qw0��3J��M�������]��v�B�ޞ��j��	O�����E/���G[����Zk'{��O,"E�����T�m�l~�(�*���2��u�+�~���$}r��(�/�>�m�a_pg'u_� ���ZB,�d��u�yv��L��ܑ�Uv F'�,�>����4���W3݀��'D�Pu.il��t�Q��sj���lʸ�,l��B���!�(�d�e���#�GT͉ڹ'�Tcx�"�������`C�1�H��X�S 5�� ��9�����H�i���y���R w�qsoK)4k����o�M�T�'��Y�ߗ�.�ؽ3�S�8F�U���d�w}#�,.ur�-p�n��}'8=���+���	���	���t���,-ު���^�ߣ�+_�_���1s��W-�;j\g��C96�.C�>��x���ݰN�-��5��X�y���2�8�J�Ak�BЖ�T	
�#ci�:4d(<�&Ӑ+��߻��ͫ�VK��"�J�s�n��i��2~�x��W{tb����z��XL�2�\���d9�
dT)�簎�����s@�����N#$t[�
"�I.�YB�[?��{�'o���҈9�UT���$���U�mb��:��
�K��0��n�����q�9���L�Y��9�:���H\#�ٶ^����b>\Ľ[vV'l�A��2c�].�v���8�����*���6�� Ѥg��^:p�H&lO2 Ķ��gޱ����~�*P�^�ѻ$�3��̤i�]1T�G��az"���(?gJ}�Ц���H'��8G��,V������k4lPa/���o�*{���;=Sw�g���鿣���<7��8��^&�ͫ�&��͠�D�=�i�� 9G��a��լ5�g^g�z&s���:v���!q�Byt1�N
�0	�QZJw6_:�M��EG�;5'٨��`��v� U�g�ǚ�%w�e�m�����/�K6	�P,����kШqM���e�x��5�l�2�.��N������5�Kfƶ��ض�pɆXA�r�g��N��:�ŏ��N)�=J�W���<l\�M��?]VV�0�6ɀ��/oHD���qK��W
�A^�&_�H��*�D�}hʷ�ۮ��s(%6�Ø+�bKn{t����J��jPZ�sg���?�%�9�e&q�0��%�uZ�R�KL�J�[<֯1�f����}�W��L1�n�l��9�j~�'d�u�oIiS@�v�G*VWnm�\` �u߅�$�}��0To���S��g�Y�	r�U�u�k���6j�s��ˤ�X��7ds�c�G)f�T����w���nZ�P�kZ�˱���?�1c��_�^�7IQ-�(~]U%Z6�IA�yr�H̪�Z������NN�1{��a���W�������Ir'QO�����ze�L��r�&�+�;�n}������n����d[��9by�����%��'TU�5��x���'��h�X�`}5���,  <]j/�`�0��&y����]k���@Pa,q�������]�� ˈZkhV�MW1+B�R�y5��L��a�X"��c�Z�y�kQ,��칍�x���\��x�R�9�D	S֒�*z�P~��)K��Id�y�q"�**��5$YPY3Sꎪ���xld���Ɵ��
�������x���U���r~�s��e�T��i+�D�$�H�^�A�> �Q, e,$�W�6_�Q�ef��2�6Bq�L��jތ{��j���*�Q�u.q��ʫ�,�է�AŢ�;�3X�n����֔)It�$c�+�V�� ��I�m�hE���^��&��;~W ��|F����q�F���|���R*Z�D���e�<�S�M��Ƨg�)��;��t�59��6W�eϲ�}�;k}k� x��+��e6���>�<��6��C\��׹�N���{�Sw9t���G \�����;8]B:��d�p�[g8j��c�X\Pw���U/ӻ*4��Q+���-/�vWV��A�f����1��!�<i�'������wuQ�Ԩ�SXqSH-�Ho����{b&ʐ�ח~��c=ZD���6B�Ǌ�yi��6ٚ�j	T<�h�y0
5�;Z�� �6s�O���D�v��v}����:�{�)_6CU$1�J�=Ac̆V^�����������~s�߰g�vOLj��U�_4B�J�5U���̆�0�ҶW9+������s�r/�P&�t�'��_�/�\f�=0�"�7T~��v�_캼Y\=�a���}����XgA�k�	��S�*J�y�k;�������n�d�A��Bj-��˥� �@�� j!w7!�����#K�Zؘg(<�)u��v�׊�X�b�*���ȋǟѪ��|{�[�7�)���E�zw�>��hi�-��6�߁O�|i�:%����K��Ya��8�yG���!2*�M.,�r�6��E���긫�g��(��;��4�ǁ��5U����t@�*��R��Ո���X^�e���6�����=�>F0����u����x��a �<%��&eXB�����6R�-�e��0O;p�hف�E��A�ol�J�����_�;�q�(��M�M� ��]�%E(J]�y�h`�V�R%x?sV��(踉���G�:'Jux��'�)�\6�1����Ț�I3d�	ʁ쏥]���������Zd���P��oUN�lHO̪�pf�2��u�)ڹJ +��P�x2�/8�'��5ٴK��rD�9D��L�֓��I@��29���<D�����P�o��k-<a������#�WL����]��2hr�2e���RM��|W`�� IV;,� ������\H "��rp9eM}��c� k]�,��ږ,C[��v��b�mœ�Yb�\��
>��*0�X���a�<�&G�n��%O��t�=ڬHh��ӗzA����'=����
���(�����Q#چ��@�Ԅ�}F�򢅭t��K�f����W�9�ƹ���c�Y��E(��"���z��?w	0�g!l �
�,�Y�{}��0����Է1X��ȽZ�'��zvb��s4@[�����y���z6�:�
?e�$��2��r��� &�y��g�o��Z�(2��U&�ɢN�� $�,D���b۷�#v�߇���(,��)`���s��u�q��	h��IW�%�, ��F�^_���SR��mP��cY�5�-�kN�}k�ѓ0tO�$�a)��c�A_i0�`R�7�:�s�(��� TG3�;z��澵�Q�?ۤWn�`(�_�b!�
X
���=e�R�c�(�5w`6�:���S�.�alcr��4� EG�Ԁ[�Rt>�Y�3��ʄyGǳ�{ˑ_2І��֍`�Ջb;�=�݃r���E�݋�1��m��'����1��r���D�7Qk:��D�}��}X�_emÎ�±�\8E���?Ѻ�Z�9&̷�͝X�Y< k�˕��n�r�`y���C�%�m��K�и� �Q���O��A:-5K����T�EMt=�k�O�+�Y�'�QG=䢈rK,��S&�t�9zz]?��6��?�A���i/�����q�Ʃ��X�z&ϱP���,�'}F��-2� ��};Ls�hce������������g6�T�@F�ݒh���au�dň�dG�֐�΢P�oG�H^-���7@~�(�'�m���B��(��7�/;W8o3����E'�w�M�CZ�x{�'�ȕ���59�+]tFO/֛�(H�K8o�y�xk��omNŵ"'@�ř̓�k�R4��� ��s�;���R�S�֪���S���s!F��
�:���yQ�Ny`pW�7w5/Ɗ������c�v�J7�p�Ⱦ����Ok� ͖�7~D���@�թ��p#���7�4����F�V*����8�L��zʑg--��.�[��q���SA��p�Ы�Nsd�0�VW1¯�35�9"bՠ�8c=�x���g����mՏ�Dc�f��xg�o���s�V
E�4��n<��{��ɵDkS�N-n����1@�t��*o�6�4{�1��"��Z{6
���_�A��SOE�K��.V�,�;�b4_���\a��>��/,>[<2Ȱŵu���	�3�P�ZomH�a3��N/��` [�����8>����ۦ�\��=�B|1��c
B>�Ń� Ia�����U���M�f|��n�+Gps*lX���"{��0�+96����5�3�Kd�vB��H�f�95������&/�^d��dDn�(y�{u��X��6(%�9��S�]�lhy��<UW�{~�.����$�xk���y�[V�ș�z���Օb��3#'�?����=�l��O�O�X�TFޓv.X�_%&��ƥ@s�8�u�{S������Ν�o�D���*���H���d��J��}�P�?�W��[��g�V��Ϋx�bv~���c�����u�@�"T�)(�=�!I�&��_U��!d8l��j�O��{�c���4��Cze�����)H�,�����-�|TI�=T���o�rbi+Xh��,�@��	�B�n�N�º/kw~4l�a�z����(�4~Lͤ#7����#��"/pt�S3��91}b1�D��
b�;F���&��k#�j������j���E����uT�.c��_��ե��������hc���3����<
���L�ڃ\`�'����ol�=�+VR��TU~xP'*X�[ר��.�ü]8�X2Y��A��so�����{�Q��+w���'���!Ni���,|�G�7D�C��`R�-c��οS����}�G䫥Z/9nz�=�u"�bo����h�ó�O�{�ls7背�OZy�����Ȣ�xR�!�v^5n,�����&��
}�� ��s�̎2�*f���W�x�yN��b4+���u�T6��1��,?2���]r�|�ͷE6ʀt�]��S\�q�#�VˠF����S|���`�D8G��[�k�R@�Z�p�wߖo�A^"�#T�����>����S�m�<��c��i�iG7����H�!xg��+�yq�a�r���:�y�E�EG���z]9|����s�^>�5n>'������D���%j��A.� Q��[�ON�,�Kb�k1m�){J�����K�0�e�_���hT��������A^��nNy�;���'�;�
QE�K,H<��M�*3`����0��-d9��q�r5���y46	�{�}Ŧ��M'��l���ОX�m�a�&�r�+��1�{�"m���}��m��e#^���.�]�	@��D����K��$�x�1�4�H��(g��rE��L�6�s�lV��(Gx�\	|K�s��|eI�u G9E����Fmk��q��I��bR5�X�_+�o�`��4����aZ�����{l�ab=��uj�T�D��oO򿥊}X�-HXQ�3[���h���2�p�F����E#�"|�><�p/��li��5k~|}�L���sͩ���0ْ�%k�p��Z$�+�UR"��6si��۽�
�����k^�	up�[��?E���NS��{�ޝ:B��K�+��ӽ�_�����;����%R>�L�A���B��ܾ�d%�P5�sp�!�slVxFV��,��o��P��ec�Դ�����^;%{r�1:�ʮrQ.B����j�^f#`/����O�s���V����y�'C~�q�QX�R-%����Ѩ��`c�%ÕB�7ƛ@�4φ`�XXn����
��Կ�2X��DCچ u%����óp/�-�=�q|z��6��=�AA��!Q�q�3�w�b	�-�(OE��R������:h�S=g7��\WO��~*0=�,؍;�I�{A�EXW[g��>Xq#:y�$�.��:J��&�#'N��]�Z*�7b��-n$��d�d�OJ���V{�"�@Դ�u>,��RC>���W��y�|{MG��Y5�
���v�s�y����\��3|}qb0-ʄ������������z�R&����I�x���գ,Bw#[O詾���03�Gp�0.<����Dp�z
�
̌�b�V����Zw��W �$�|��c-��K�'��י;A�b�����GHz�V��O��exJ�����qK|��)�99?)��㑑pQ�E��axH���B�a=01�~=�_7���Ũ���P��3�9q~^�.��a��+(Tx�Y��JK4u�O��h�	�̋�ܮ��U�Vx�`�h1/}̅&� I����-�Թ�j[3qn���XH,uvӝW/��TqT�Ya�o�D��K�PJ�]7��:I�����bn�� �	��rL���.8��X53���~"������0p������UH�Y�M����?kj?���}��w��O�*��\D�ުAUߤP��3/bm���a�����?�O� �_K�k����Z�f�����6SY:07�3	��t��-d�ԝ(^��'σ�2�����d�p�� �"�&�͔.���3%�ǐ��q�q�z[࿧��+W;P��rI�{}ʠ���@Ņ�o��mi7�۔�r�|XW�E�Թ��mP����)�?�f;���`�x�5p�=>����Lj�i�xh��.��ѬeD��E��c|��.=U#�ľ�������D-�n ���3R�+�B� |��p��Nkd�G���B������#c�c0�Z���m�.����<^���߹�q�¤�M���V�����q<mA�~�eO�׍9zE���%�I��$c��\Z������J�j���,�:P�ǆ��`u��T"	����hx/��އ�`�/�SxF·g�?��TZ���]ѡ�x vԑa���`������Åɿ���*�[�R!�JA��ڑ���!$�F�:�2	�Co]���*����:P���6q0����J�+���d�#֕�&�*��u�Ow�)դK-s���u�[�6�}P#=�V���v�8h>zڲ��3n����������QVY�M)�+�C��\�~��0wYl���5�yJ���07;���\����9{�Ӈ$Xذq<�5���Oг��ι�z�����j�o҄0�Ϭ��?c�H8׷�T���l��̬h����$է��'o��3�n�t�~n�<ֵD�zS�P8 ӝ�\�����,���U��mQ�{v�9��G�{�X���ƍ.��4���%q�����3��JQ��=�zaڴ�M�Tf�3S�z���Qߖs��p].Rŝ�]��]ZZ-��JL��V#mJm���_���?e�z��x��Nn�S�ɏz�j;��#�;b��! Jl���-�'���%��V�ek���>�D���f��
�`�h�;k�
�Q������&��s{v"�$�PWV4����s���è��j#�� �c׻�ӟ: �\2to��V��T�@Kq�����}�/؞��@�>��[g��EeD�z{�am���U��u[��h^h���PB��I�e���a��JJ�w^���Ҷ���sp~�$*gޥ��^���w5��:@��gA�"�\����~}�{���Q�zo���I�Ge� �wf���W`�S:Y$�x�?sLϊV{a��G��.f���߲���,��[��s��#+�XT���rv� "��d�I�E6�s�S���s�Zi8����4N���3p<�HJ�Ե�p�t�����@��7�;�Y�C[�'Aj���i5���.�x�+G̿I�.��]��_�*�<!��-���9A��]/��]�L��?p�j"����"�s��FYW7���]�1ok����f_��u��G�)�=7"��R�@�Ы��28e��C!�2A
L1��ɕ���[�id�HK�&`,[��M�yg66��=q���F�b����(�j�D�}��=٫�����c�	z���&�9nR����q�i�Z+����ʩ]��+�D���h\�.��9���,�N[����H)'��\�v��M.����g��>?n�M!qB�hy�Ԛg`59��?�j�x��4E����*b�Zj�ș&�*��N�[��B�G!�L��;��:H�r�w#��|�nӻQ��$�c���J�))ԍ�jy�sG�\�JTn-u��j���R?�v���{a�}�?��Yg�y�݋uJx�rI�]���ke��`>d�;�-���F�`�Q{���|��?C�X��k�5�{��@D�;��/�^)r&���ݧ�,ᜅXv�L�H>�/L�ժK#���w�ɔµ��N�߱� ����?������@|�RDK*��d���#&G�Z2��k�Q�H���v����&�/`��S�+��;����ړ+P��[t.�"�#.�I<")�oB������8��5u��T7�Lr�JsJ�h�N��h|���N�c�0�k*��0@�/�!���g�p2�V���ټ=����G돽^ Z1۽�뻔w�@_b-�~���0���!泃����!����>���L�p�pl)XvM�b2���J���l��i��g|h��A*�9��5u�@;gy�v�%T��Yi��;J����c��oQ3���,�6)c�ۜ:r7Ml�Y�mG��H�
,�'�!﮾�kW&�?q���;6��)ţ^�:���`*VⰎ�qV�a���"2%G�/d|`7U��m	�<�����Q��<>�C:I�j:����(9�zz�#��q�S�k�����^��w[�d}�W�op69&����_��e7����a�5S+����s���\��U���S�x�	7�Y���)@����Z��6��_��<�'� �-]�J��$?�%�~ON�*�5/pVz���L��c*׵�o���w��h�7��Ƿ�f�� jų�I��s�5:��>=���s��:� 3���%pK�DDi�#��E�A�NBk��ܰ!�g�C#
>3}_�p��s�i����g9W�`D��#�嫂�%�{U�(k���<��>WNF�io�_x�j��mv�c���� ��Bi�	��DY��
e-����'B*Q���Ă�`�ߝ�q�7�8eGƥ��:��msMex����\�����K(F*�L4v慑�b��A�̱\M<�~$���J����Fii���H`��;�մ���Zq�C��2T�ĭ� V5a
���	/᫽����	�h�,USY��L|���>(0�b���F����w ��D�E�m��n_>�+���XNޠg�v�븋Wc�@��L���|��'�+��aH���E�����F0[
�����f'Eq�id��7�����x�M��Z����6.��cA��ІLS *Q"��z��+�v5�'t��I�H��������=S~o���j�C����Q!��\"^&ߛN�ʑ7ەz/9'��o�W���8������Z��n^b)m�U�b�O^��9�h��Up��
u�c�����]o�^�m����9I&��	\�D�����T\��p��FK�w�ڋvl�͢u��-^~+i�iNL���l����D�X�-,��#N���NI�rCRfia�A_� ��b>1LܬF)j���F��B:�.k�M|C!�>�ߚݻk�%����裴�~�0hm�q�EM�!F�	�r�!�D��� z��9܋�ȹc�5��^<K1��+���מi�n��:a��uծ�m�F�,I�uъ���E.� �'��n���c�ba~��H).�o�XA�Rn��mct�R�k�u�S�r.�)����[^s?c~�  ���x�!~j0ϑp�7]����и�lzXDA��m��ԚE+�p�r��t��	���Cו�w�54s�;�NΏ��������(c�������q�E���Z���G�������=�LQFV��r����?[�ֱl� ,����$����i��~�l���&hv�rb�kok.��OP�B�i󬳡�J�R��H����.[/,�ş\4�S��j���+b�1a^a)�S��R�1�T3/�����),�euUQ~UY4�=���o��w�>i�!6d4�S8S� ���⠽c�8na�޴?#�:b����������A�0�8-Iڞv��3O�#@�" ��VF����@��
�Mu�o�6�lVCO�t`�;����o��;91>�|'�;���6��r7÷���s���$�/�`cp�l�	")�Q�z��(;8^�@�N��s1-)UXd7����Y�:���������;�i��i{���|r���6!�l�>F���tc��!�3�C�*����^��u�f-�M�͛���)��'l'�Kw��2��P���$y�pfC�\���{;�z-S��(m��[]�Nʥ��\�������5Ha��	qƖ�j���ݩlJ�8L�. >�C6�4�?d���E�$d�]��FO�`��#�^�:����'$�9�qD8
E�&�����c�i��c����U,;�ܘ����Ǵ	B�~M5��o���H=q�6J�SB�����]���E�n&�0�{�񨁶��,�w:8�j	J8$�������T�8���%Ƿs�a(:R@�=�8:�b�O�:�\��R	�5����Y��~ZI�`Gr���.&Pz�b���[|n�$��Z%|��^@?"�z���+�y\�85 �1�&�Y��2���+U�:�}WHnr��JD���k����`����]�GI}1�t�4�%��ӫ>���~��ZK�z�a#M܋�U@=�"�=(�J{Z,:j.��n1'�l�䦻&�Me�M�-0ڪ�YF��p�ሑSR�c��RL�a�h�";5�-����'����.��- �(R�@@���W�Y	�VTش���O��g���4�9�j׿eY�� �#���Ƌ�?((�(gvp�r<v��Ma/�UT�d�1(oE{��v����XP �	��Ze�����5ED�\�x��Z����,C�������et�?c>A3v���8���w����nd[�U\�/�ު�:���=u{�]�Z�L�  TmԱ�\����ǌ�j�1�K �Ҟ��W��vL��0��ÓLj�E�#����!A`iL�^���ɕ'�gȇ�4���(�-N�}O6W� ����LG~�/!��`�<����Oe�yI���,��o:�k�\��aPK�&t�A�#� t1 ��糇�2��2�!��S���K�
�u�Lx/Yu�I��j���B���a$���,��I����:��L`%�}3�s�گa!Ⱥ'8�ߔY����~w.�j0B�ȭ��z���K�C����r��n&�K��fO��׾�x$/�?$��w#�+�w#�C;�=26����7�V=JAu&8s���,[�� Vm�e�,<I���!��\�vΘ�D�������=����F�nl��[5��}����,�H����6�^�1�"�>V�{Ӻ���e��l
�~�	Cj��ե��������w��o���ӹB��v>!�w$&s�=e�f��j ŕ���e���`/�6gI�Y�y�%�/ ��FD�u8z��/5v�|U�����WᣇU�Kz=B�N�/���&����į-�u۵�����;Z���E�}����Q��$qI�0���:�u�Ò�����/��	�Y���(��e��-Tpa��5����,��� a߀��������K�"�r �G3�3Zac�-�C�	C\�p����W��c��P8yǀ���}��Pl��̲u[�8=@�x����ϑ���:g��g�*�q`,-x;`��s����O:�(��E�I�m��S��QHd��, ��osܣo���_�<a��D5�\�i7�W��?1azy�h����vLQ�~�/�>�J�΂���W�-�ZQ�ڡV�ay*�)���^�!���Y�I� �y�e���G����W��W^.�h ����[��a\���Ǳ�b�q���P�;Kaސ��h�D�jx��R�I�<��1����g�BJi�կ˷�cse�v��#�u�]��ք)|�1 �OV�c���[��P�-�@��� O�_����$َ�$���Q�~f����S##1R-�֒Z5�(7�svZ�{�j�E)�M�W糄e�s����,!d�)��G#��!Ank���Z��\Q)��{ D����ޠ�ي}C���Ɖ��l{��)pȜ�� \�@�X�G�@"?50��s��q6�h���!GW�ޚ���e��vEB\�*�5n��F�{tR<�]a�M���A+�U Ԡr��������(�;h4��������
-�?��=@4a� ?��5���32v�	���8��Ǳ2 !��8�׸Z�B��:ԏ�;�4��UA�z��E���%�w��'G�V�ז�٦�w-j��<����@[�'*@�9�d�flg�ə��	�n��续�����8�#���	�:��ѫ����X�����h@���#���4-hJ�s��;��k֫���$�%�%�y����vs/�R')��!��*5�Na�0*qM0��E19[�I�4M�NR����L<q�iX�2֮��:�ϊ��I[ω_Ź�C^Q�N*ҫ�P�R$�,��(��|�Ȳ���<�h���::�F8�wae��BBy�e��wU�an�3�GU�&�q��g�R����I	�`���_C����mzޫ��:���F�vg�2��`�Z�s�u��z�����P��F�OfH�$g����(?��"��v[kX� �{��51�Z���JS�'x8�\O�)~&h;3�?�ҡI)?+�q֢C���sKq�EM��ud42�F�7�7)�=�M]�F���I�[�t���@�k�+ϣ�
5�͡W�����>�����#8#��Pp>���҃&˷\l/Y��(bot�i������XoV޹*+�)�2��h�;	֝A9��OnNr�Q+ �m_��}#�������:�-~��G�?����W����#C�!��H��,�=�r�+�]�,�ۥ��a\V(��g�x�2�(�NuE�ј��q�Q�sQM�6���KS��H�W#*�$f�>C�m�$ʚ��g���K����j</G�w�]B�@+�,�P#�A�I�h���Q�J�-&h�7���j�d�2����q��I{�3R�J��i�e�y��N�
��H�E�1��|Ų����V8y�t��'����0�x�*-��L�������:`c�������b��k}��2��\qp���&�Xξ�>܎�`�M��!���Lʢ��LH����&  T��
��z��C)��t������J�2j¡�Uk��)׶H�ϪE�|3���86��bi!��E>�H�kaU��ǢS��U�&<��ƻ#���<���:r5�K�[��IA�`�Ǽ<��D��v�Y�$���t9V��o���`����:H�Ɩ��$�O���YͶ�X�;F_2&h2��!���)]�$m&\F;'������=����$�A���+죺���YuV��
��`��9W�J���@�l��%���sg��F��ǖvw<��5)%��<3��zH���P>��mR�2pr�v?����K���TO����LO�:�����Α�:����ں��2�Ie��~��Wť�Uꧩ9Z�'�w����l�Vt�/xC>�Ǥ60���,�[�s�W��~>l�nWC�)0���׉�E���ͭ<1�Bp؇��E�(��2V���&���q�W��\)���%�Q64W4.����S� E��<���:pz�nSQ���3�vH0m�3SD C����,h���8Mi��ʩ�m���&�՘�����e�f�Y���أ��8�w?F���t���6>o#�*��YL��|E7=��uÎ����ʯ"��F4ֳX�O��q�j��#=�e����Y۵2ma�Y�ٛ3SbA�p!��҃���,�<��B�hE9'����cSc ��`�J�^ܥ�$���m��$�5(6f~T�a2�|:I�t񘈳$a�����"�S%�|<<�/]�9f1:�d�*��b@z�ë�)�Xw���#4᡺әL��O�� {����L�1�?*)��	���!H�@�`�RSΦ.�h��t�o�����߭��;�Ż("�V/ZWt�� Du�``��z^�̞�y\m���� t%�.�]z�߯����sx@*g�z��M�[v������b s� N��/��^�նn�;�C Rܚ�|Ln�vڣ�~�4I�gC�5�Ƣ[��F�&��K�x���&e ;��������e������-2��M՘FZ+���EU�Ft�^���6��TZ�g���@6�ط7�&��IX`I���=|H�0M\�ތ�[�
A�"�% �p�.RX:-�g~��NQ ��� d*�Jm�x�� �6�$��9�r�峺����R��gד�v�&	��Gz<�We��Z` ���s�CpC ׀׎�yHP��@ͤE[�� dG)�}�^�(ͫ����.Y]�wM-���!�"��K�킾%�B��+��p����;��J��r�5Ǽ�w�w�i��'a�����[�X�z"bg/=q�˯(P;�m��p��[=[��X7quu��?[�&���i5�`t�N\�!�5��X�>ґK!���Ħ�(BodOF~ƵZB!;�ΈC7���_%���:���B�ֳ"#� :c�h��2KlY|�*)���j�����Cߓ��1�S�fޒI��W�V�@��4~�����v,D�8G?�=�?}[�C�j��w����A���(���};�/�:��a��T��2UiF�٬!���w��>O�~ �xځ���/߿�7m��U�
�Ϊ��C�GU�'�2t����e��QaA��rL��,kU���s Y��P]�>��=��!oP�~�pˉ�{U2:��RlB�՗��^.�8�8؁Դ����*���F�h�,�8����D`lr�ش���f>H)h�2��K�>�x`�� j�o����|7��1��T|d�?A���S�;�/%�c�[��
���7~L���Zk{jm��	UA�N�U���|���2"R�}if:��Iwq����R�z/�3@��la!'+��£�5�꿏8�`���A��i"m�ћ[��:J_�o���%��� �.E-!y�滋�r�l�׻�̦6S�)9F��3�q9��~c6B��o2p+/+;��,Ԙ��P�fS����4Z? e:ԑ-�3��V����+�i`�����g0/Uu�k>�u3���76Q�Y�ya������B�1F�8\�2���5�!:y���z�X����Ҟ��:��Kr~-)�r���x>�_o�/����V(�`�D�z^���&��ʴ�[~$1��B���d�˰�v�:j����?�=l϶������x6�=�o��r$1������3�s�htD�����fi��S� �3i>!>���f����h�W�� o]O�Y�a�<B[��~��#5f��n,�D<;b�N8,5@��P��!a<�:Lȇ�i�s�lr�fZ$�i䦷�AfKL�)��j��Z�>����/v���4���-`�\��u��"�R��2� ��]=�ſb�`@ΣR�3�ۤˇD�<���5�L�[T$^�v�.���G���E��<8I�eX}�hMt�m�U4�W�Ā�1�:���6_��T��k�ٚ2�J!���#I>���ؕ���Q��["�9W�����%��Y�z�g�1��Um�����If�ʜ�9wq��*�^�).!mi�A�c�=���J�z.��_!S����χ��o�Z�~��S�� ۋ{c%��a4d@����;�M(����}�B6!3mڮ%���K�qPD���*]Ƿ���h*��.7����W�	x��t먪�#�N!v	|\�>�^��Uw(���I���^���Z9%����1]��YÙx��4*,������
3���0� %�o�z���Z�)j�fH�E���3RqY"=��]l\��L��"):����f�Ld��6��*��/bt�N�
�m ��!ߦ6���N��F�Z�L�>�3VA���]�*Zd��2���:A���1Ƌ��nk�Fj����1�,��s���[��L��B�����}cL�^'_9���1�Y�I̬?r�M�9E ,�r�"xA�V��EEB�E'�����Ȥ4��j�T!��
���
�� �d��Z�S�1'�����,^;�f�L[[������-9H1�\O�9K�eTW�j���/���G�jLΚ�3����j��N\(�z�lbC�tI&�@sx��O��f�!l��n�*�����b����1�_iÉ���� �?��C��2L������v�G!����f&<{"�:j�������E@����m�#:/�s����]��=(�a��8�z7c�����*}o��H��ݩT�7��m��J��~ю�����^�S�����,�����.��lW���NN�`P����Z�JY05ӭ�J�Z$P�)֜R�9r|Ul��,�D��hy�	����E5�+�*��x��y�_�@���^�7���\I0M�MX�qIy�S�c+Q���(�Hp'?� �.ہ�#<|h�e�O�%li 3I��4���F��Բ�'-ޫ�M@f�ʖ��3O�wq�g�x$�3;K���m���`�Α�L\O%�f�%l΄w
��1�v���'�B���:�k�͊�Y]s\�}]%Y�1��y��^vG �p�C9I�iqֳ�,0/�Z3���ƛW��/�Z՘-Ϛ���/�>���;
��qh{�5M�v5�Nڠ�=����9y���������B`�D�������qcr�������8��J k�ǔB��[��Ȧ��]5�9�/�^�ӵ�	���z�BEG��Ob#:�<�_��XV��W,CIr6������pM;����j����ud����l�0��Mc/�}��Ѿ�f�0�P{t���T�Μ����!S��ܨ��/mR�Qt�%�y�����o,\���.ҙ<A�?�F=��#�EQ��������4j�!�G�=��`���9��W�1̹�=j�8C��0EV]�%c�5G�b>&�w�'������y n`�M��[~�2 �@}�
��xZ8m�����_����F4E�]��ҫ�+�����X���`%w6�w�Q��g0���۵@4������@`��M��GxH,�w�jrSțD�l�^7��*gr�Bwج�U��S��妡�I[�C�B*O��
�488M���s�,�]�Rŕ�K<�v���%�w����q��0}��	ɽq̜��ub]�F�ߙ��z�-oV0�\5�qt�^���m����$ {�?�5h� \�����,��Tg��i���n��N<DNIzN}����b�t4�\�4�.��1�E��UBt�Z�q:VX�-�tx�T+4�D���آDϊ4i�H,9�0�L��7@U�Tެ�ɊT�5Z�(`����ćv`�шE#+�����d��"���?���A��>?%KHW�zIe�{�G�B��d�;����ayg�͟�r&z���=BïljZ�_9�7&��r�H.�`I��_�#'��TBW��Z���h'�?H�P�C�j�v��%���5KA�[Hlba8a��+�֓ ��E���2�$d�e<�U��k�����C�By�˅W�Z�~B��Cpzu�_���am�Eb��ݫ@��[S�[�0����JX������v��|
�d�mgjh,��������k����0$L��VLp[}�cC�oD�7�i�4\� *z�u�ؓ���"�0D�?N�%_ܦpe�z��(Ԕ�ۇ�v�E�G�����;�;��d�҂�,G��P����	��J�PN��sN�`���%�듻b:e, H#�P[�4�u��S��"cʂ8���PE�ph�Q�|���f��G��e������^��z{AǗ�aeɱ�V�k�#u�_\���2vĥ#j}��9��u%<[ �p$ f���d����yv�L���9\0���d�֡���hfy��{�����$͖��t�f/"�iW�K�dƵ��˾��ݒmL|pԦU�/a����|�iAF��9禲�F���5��pj�ٸ��F�B�c�n�R���ȩ��^�'�Mf�"�NO(h�@�di���`x3��ǁx0��b��2�v���2�,F����d��i���pf��c�W}����!-a��z�^y�o��/H7�b-�w�ڻ<�P->��}�z�#�T�ց�[Ps�7o
�e�v�	�a�.-�IQB(_n=��A^=
�<��sw[�½�ޙӥ����v�)�0��T3��ssx���&^`G���<�l��#(�7���MˀmuQR����sa�"�*�Ԛ��y�{�#w��1!�<��P0t�ά���؏&�V_�?�/��:����A(}@
z�GV[�g&�j���' f-]�Y�9h��'�}����+h�{�JԱ���h5 �B�Ͳ{�HF"j���<Q�*�2��e+��>��=�(�����cI8�(�'�z�����I��G$ۊ�<�9ByS�Q�|�F��T)��Ȭ�g�_|�ѱ�~�G�)H��+��ӡ.P"�l`����YMU�g��-��K��n���RC��F�f�u3kO�;���Z���GT�f�2�J������ej}�1��d{��|�hJ);�!���z���c�Z6�c�GnIni�MO��_ޑ|��ٺ��ٙ��������[�	�=�������.�2��%���$�3I�Y�욫�TQ�~�X"�U0P߭�x��[U<ڦ��:���f�=�O ��5��88�a(rEh7l2�$�����T`��k��8�N���]e}�پ���&;m�EP�Q�?�"�c�z�.>�H���U��O���G Q����6_��(%K"x��=�;�lecij�j)����h���1TY�(��q��I�;��b��u[�S�-��A���A�#AD��ٓ�������r0�J�o������d�'xo�1#?u���Iv������xTa�a;iS֩f:{x6�_��n,q��@V}La���c���æϦ4���zC�l �������i�@Ҏ������ %S8�H��w����Մ�q܉��sJJ�_�b ~��^��粣��o�����C���x�eqm���ICa�S	������K�$&|���4,�g7���J�S����m�!v�#���qs1I��i�~D�t��t����i���߼ȼ
�R���"����_��lf�y�	#ȉ�2_<r{�n�[Y-��dq��M��`K�����Ln��@щ\c�'�g�p�����3x>,� �GѶ�{F����O���2F�hkzM/v� ��O��:~n)ޛh��ND0=|�&Ql�#�G�C%��_��uv��_h�X����I[):A�[�����+�t�E�T�6��4{����������u��.�Vuh-V��~4 ��?1�6��ҎQ��c'��䤫|_�X)+.܍~�?���vh��vđ+]� k6���t�=8����`���t�1�VG�y���H��Flp��sV�kot7�Bh��X��a9+�jx�����$�:5u�>L�I8���0D�"�X|5"(y��Ȣ�e+��c���b�n��ŉ�]���RE�5�� �BB����֜��ۮ<1���A���#��� �E[�6Ӂa�{�A�Vս����'f��!v�?�O�lr��`�$/k|tS?e��hzJ�����:<.�x�8�D+�$���g����O�L�.�,䡂o��K�=̦"�ڢa\T.�p����C\���O��񊚶{˶/)ZHL��D��qa#Ⰸp Q�R:Ȇ�Q
��9N.'L�-���z͘Q�r94����ݨ��
x�#����q�+�=�YnM�@���R3 s~k�Ba|�$��|B&��!��qȊ�H׈k[z��7"A\)��?��2S��k��8[�,�I�㊉)�#���0�F���������) ��.N@�)��ud#5�U��,�t�6����C�։�A�swp�r(��E��CC�%>˹�;hnӵ~��G򂂒��6*�YNB>,�䢀윹6+M0�H0W��`%#�b��c(dޞ��F;
G����ó����c�c���i�a䄍�S
O�P9/��o*bԯ����a��l�I����!&�TUd�OA].`!Q�X�w�2�x��ivK<�G�sW�[9������7��/�v-��PxG `?y�v�����.�VaІ0�hkr�\<�/�G����Ҁ���Z�=�M���|��(4k*&��6���oef�*ѧ����e ǶG�`1ؐ��@��̳!�0E�6���:��J��$�O1�g]!��X�^3���YD:n��7�_��?U�R���� ?��S�I�"5Lf3�"�6���֪[��y�/�<��O�6����T,�w��C���g�),�����t���x�c'4S)3�]�N����%K������-D��6;^�Q���/I����f5Hl.t�A�X��8����;q��zK�]���-�;��VU]�[��`���jL�o�P�,���85�0p�fOZ��V���A��rX��.�ἁ������~��6NR��z�W�l=$��y�� ��CL���s6p��@m�^/l��o���s��&�MCu��C���Рǋ7T&��W��d���C?1�����u�H�=�o�Q��cN�E/�˷���V-�	cTN���n���*X�D+`N��y=�P��*�:'��o<,_أ�ښ�q�����d�A���] W2|Lqq[�a9���[1�&��	(���Ţ]lp0����.=��ߤ@P8bg� d�m�Gz�^��/w,�k�6�ZIm:�����L�x ���>�1n���ZH�xkh���]K'��g�4T�L$$i���+�+�!�
��w�ӥ�T���s]���;LQט9|�ŗSq83���uX�hT��td�V�>4#��/�/H� \��T4 �M�1s{�O� �%���
1��+:�+:�%t��+���<4���4��*4�+��=ʢe���4�����*4�󠐎l�����S�:����3�gB){�*{1W�=?�8�@���
JV`�>k�PY��c�������8���� ��)��S�GO��R:���{��=��f��wV�����T�~gXw"���6<5�y3��QT`ޒfA�0;��Z�_�$iB�EH�u��a4Y��眛줾�A��t_f����_�{��OE�칂zp
�;��\��W=x����[���5�ɠLa�ap��l��>��y�m���wX�l��s\Z&���:�I�QG��]0&�ibI"�[a�������]iFs������)�#�ʢF���`�����ZҨ�z��ZE���h���e18�jm�'�w�UUX�(���rI_S_M�V��`����X�@i�z�WLX��ĆQ]�)���[K�������AI�˧��$0\��\GYɿ�!�]+ǎu��Ċu�4nz���@,U5D��o�eG�.7����1��d���>��a��9Cn�r�s0���#O �>�W߇A;y8��]8�o����n��[���r�
���ӺW�1ry���o�Y��.�
ޤaJ2J�OK��%cX�CMp*��3��ߋi�."�d�2]nhh�n���@[bn$"�@P��f�'�_���)� ތ �5TP�Z��|@���d7W�e�������
�E����\, Jz�]��;����'j���$b�f?�ڮ3_�'k��;M�F�� e�4VV�������Jx)}���T͸���})
��".���z\Ռ�j ��!��g���m���	I�x���,�a��\=;�G|J�(-����3d��򧔘��T2��턘(Mi'�4�Pz� }9�A<lP&�*� '��p>)<�SDݺM�So��;սv��[DQ8�'��M^���v��\�T�T��Ho�؄�L��^�_ZO�����AW�*�C:�1�N��)-M��23�//� a������yl`zb���n�2L�Qc+�+yd��Q~?�Lk;�Zr�i��K�$�9~�̾�dʣ[-.�;Q�#���R�r����{r;9,�a��I�i� ui�_���;�����6u��1>s9knmaV�?N��H�hb����!��M1�([��n\,�+���	�f"�.=���c<���v1/32zl	n��U�|���8n�F��7"���@��a<c��چZӟ*L�pkI�a�dA1�M�΁Vlz.%�r��d�Be/ʟ5l]cKS̶�R0�F�TO��N֯�]�tyM�G�f�2,�%�+ �аv���t�.RM��=�CjeA����ԋ(��K�ޟ_F��e�<��sK�.�}qǽ�k�����5����:o��T�i��i>DoA��Ĉ*9&t�p��Ϭ�D��ξ��
!�8�9���;u8ڡE�2����q�~���9^(~(��;�E�j�q�C�*��S��ft~ԯNgo�PC�M�@r-�R](��P��KG0Fsg0Q�py��r�7}�\�k?-;�{{+Q�}|��N��f�|�>b��qA��?�6�j�E}�<�"HɼY��y�����k�5g�B�*�O���L2'�>Ȳ1���)^�Na���[���Y��гzu��� %��"gK
�B�Û1��ꂛ)o�7�}Q!� O��1	�|�q
�{����Ǭy(�k����%T+�G�ݡ��@�#*fb�8n܄)��
:"W���s�{�3��
K�y�+C aڶ�"���ƣ����?GT�V��]�z��~�	a�3f����ֱ�M��Q�r����X���A�ke�'r�9����yǨ�Y|*v�̣������B1�_�5gOL'*���E|�d���_�<%i����������S_�
N�r���Բ�T�rx��s EQ#�}6�ךaU$>ة�\gS%��˜���W���ƅ�B���;+2	����8�x�?��S]����H�]}��q��#�Md��G�_�ʏ4�^`�sQ�tF���I���M�BVXb�IGyM��wV�~P�0:(Z]�ñ}��O�9 �B9����j�Gը`Nי6�"ڈ��C��py�A���a��嫰☳�/���/������X������B���pO�����9HZ~��=���Zf�Q&(%���U\�>����m�t����\�R���+��f$k7�/֠�j-4{�W���~���g�c�~���t���.|�8ڰ���U���`&>�u�_ [�>��ޝc7Ƿv�B� )��>���
����=V0���u`qp4�	��W8�f|0ҵm0.�DL�����Z��ͥ��w�w��@(^>��T���g��=��r<�O),�աK�?��ǰ��:��Ii$�(��B�~zI�˸/_HTSbd��%�ߟ�� �DnB}�J�J�?Kum����#K-��,�?�mF��lB��e]���e�K^���G���Cǈ!_�r��ݑ�{o;]�T�N'�$�S���y���]�e��|�@����-�"�~v���:����9���rT��ew�� [Y���"�ƭhy�����2�k+�Q�!bct
�6�������O�'���7�Q�'����m۳�**��P#Xνj|Z.��(��F����i����nV����LL�8{�V���نXR�¦T��CtQ���Q��aՍ� ��V�v����jb,��w�5�g��V�u��bx�w8�[� u��5�Vs�ZKq��7i"hM|>�]�O���'S4C?����$?ʿ�h��T��%�C_����}���;oE�c&�8@��,�����Q�I�5�)4nء@��K��C0T%R-C{�8nQ����q#�0���k�e"l�7��݉��x���L\�8 ���dI�e���T�%b��a��_��@N`�~��NG垜Z���J�S���ྫ5+Q��9��3�&�C�N�3�tq��&��t[�RBx�΀�x
�3�#�7��®����l���0TT�Nb�LShS�,I��'�yK���v J�SI��%0�1��V:qEf!��ǯ;�M�I�������Ԫ!0��5����l�gE�7�~��I�N���ɮ�k���㥬)���*
�n?ʣ�*+`lF n���~��y��T��Iӈz�a�X|���O
�p5
�vA*��\J�l��>�ç��9f�)e�i�l ��*��̻x  ��*P�v�f���V�b�A����(�A	��ݻ@<:�$[�XPM��)(N�ǹٶXRs��3̖���5��qQ�=@Tf���f���C�u��j�@�����
[R�)�+TY��{�D�^�^���B -��y����ud�]sѩ�i�v����z���B|h"߽�Ҕq�>�9-j]���6��I2>��]i��,�8�I���c#��Λ%�D@Ì���>�Z�h��H3��Xi&�g~tQE��2�T}��܆u����L\�R{]�}�-c����X�-��x_n�4֐nv-=%Q=��P���E�P��6zlVC9^�+(s�k�m.E�%�Xc�YI�8u�!	��N>c�<ʞ�����^au�{8G�JY�����\v����C�ʰTK��O���8�{K?�$���c~={�S�R��r-+Lk[�%>0)���aaW������]��2 r��Μ�K�WHȡ�;�]R�#i[��=�G<�WeiK�ԭx!�rD���"_%)0R���?k6d��Lf�����]!�I�t�jr�ú2h&bx5�>sU�?$mvɵ5�f:�i�\���m��V ˌ��������'�d��&\!:c]Ku��n3D�X�S4Kؓ�*�W�����'�=�ݓ��]	ػ��>R]�h�(���f��`�S��0tn/�a��4z���RV��?K������P�E�l��\6X���x�m���6EN�	�cט��l�?�RF�^q_~�P�]"�.e'���/a��=�K� �a�1;��������%j�Nn�`�$�VO,��MY���b�c��M�4���ֻ�2B�I\����Ћc۩o!�]SQX���С�}��n@K�\��E��m%�V��/�	�!���'E���w�@���e_-T� �(����S�\@��;N	�-29E4���!$���LY����[����7i��Ԃ`#������k��X��c�:���
ᒇ�����->W�f��v�MJ_+�Bܔx���y@�� \WZ��Q�U4�q��CȁZ!�����͢�=^��P�v`@�B�u4L�]���0����*=�E��Z_����}���M��Ԃ����%�>e�E� ��=�)K�'�۔� ��i،,4���hŋۧ���B䰇��8�J�y�S��i���4�����0Eg�^�-���0��Lo�.԰��.��&f�~zL��IͅuyQ\�WO�����0���wK ��ԬM�M�w�db�ʚ'*	!�!�9�e��&wy*W� �we���<J[(=o��~P��|������t[�͇uu�m(?؜����I����#c2P@���HN��TH�Y]���	1`+w3M�w��u
�#�>F��i�f�t�뒙�)P>.I	*�3����M��?�BУ����\�c��ˮ-�Z�UƢ\�@iA�"�>�u,�
|���G��Ru�1�*pT����~kw�U�.����u8�kaoMΣZ����i\�X�H��t�gWL�l�-]U2'ҿ��Z^��+޽���� bI�R5��s��-~����Cq�Nc�!h&�i%z��H ~Q��:���$��;0��]+8�X�~�.)�f��E�w�Vb�jA^b�����.�̀��͎9�E��~r˶ױ��e&�]�Ֆ�D��j����?����(艍9��s'��'8�V�h�KRwCKa�}��-��^�Dؽ�B�	�ۧ�C�D�	R�֚��ׇ�s$��DmX�E��))�W��P��u�\��.�:h��|%�	�z�4�'��'3
ȘvSS�RO ��,
��N�|�ɕ��}ˎԪm�>�24,nCwFR2�w�Z��+r����G.'�d�M�Q���jl��,��BU^�F��}	@�~��#Ν�q,����q̟�D-Ԑ�t-�k`%���k`��`j�8��ٍfѥ:��+H~�"rr�m?��9q�?�@g����[ʙ���&�[��,�O��S�Tc$<H*A!��F�v7Ob�K���<�M���~�L�I��o#��F�9`K�FՈ�]�>r�C�o����w~��e' ���FL��q����:pGE��k ��z��+�*\g��6[�Ɨo��T�:D�J�.�sD/�]=�P�KEf��lԣ45����bfh[e���>�������e�����Mo �,�e�pT9��0k{��2$��)�eveQ'U�e�A��W}�:Ӵ�ɾp�'p�G|���-��>�Y
�q�	�'ƫ�9��#Pa>.6���LT����E�B��}(ӹ�{�Y��+���
�ŊBJ�|�$LꞶ���� �W�f����J�`aVXٚ���Ŋ���Ip�&~�xM�O����c���:�X�dLNm��%���)Y�C��Q�>p�&����uyW���!7���q�N�~P!��b���i�-F��E>�����I_B�)��?Vg���T�Ŗf�<oAʸ5j��t����i�Z@���v�͵L�}�����I��6����|��n���a��$�ܵ��.ՠ�
�/DS�f���hXh>UǞ��"hIr�r�|@?X�均�Ts|r�v�finX�����%g'7��ij#���_]"�ɯ6�m����l�wN�T58�6��4#cO�	��� ���}k�-��+�
L2�	}3���a�XzD2K�h�'�� f.��9�
����|�i�n�v;��ѝ�1�ٺ�Q�"v��~]+:����TS���O.y_F̲k�S -Z,����:T�z¼��A�g�~ R���@����o�.�՜��@���*���9�����$
Ъ(H�?�}��q>1�Ю<���qU�x��)+	��ō;�c��
�2�(+���\�ǸĚe�xSTB,Q�8�r���@�ƹ��k% �%�ˮ�/DE0Wkw���N�:I��,=-n6%��� �1d�M��1��D�6�!��߱�Ζ���I�zػ��*��+&#�DW���E�:�� ��J�j_-�u��R�A���M봧=jם��w����s�7�>�(o���r�H<����Q���Փ,����I���p;��O�?3s�������L�FQ{���3�������q�޵���aq��{�7pЈ<��3�����+�.C����G�l�g:���%@ќ&z�]��U*�T��r�����1lG�4V\��c��?eC&xCf_��A���ޔ����H�Cz���Xt��ٶ^Z��?I�q�R�Q�'
joro-��+��ǫq{�u�-1�s%T�+����UY�N~�;�%�e���N�ﬗ:K�;ZS� b�f�I��\j�<dߞ6�N��j�L&-�j��~�@��������THm*(p��J�]m�_p3���_q�R���ǢX��u��~v�l#Y
,��ޑ�V: c�x`�'M/b�<�XU�f��(ж=69#�
X>j+ߔ'���#-$�wc��<������T����V
m5����MBh�CK���b?s��"GsW�̟��1|	MLi�&�IF����%�Ї����hP���E�v����V�G�(�l&�Ғ���~n���&%�4��T�k$�ǭ�A
vj�VN�� �~V�����϶�������FM�|�.�.	aϠtI�W��������hQ�>S�zk�J�Ǳ>��2c��l��Jю,�LE�R��Zؠ��Uq�-�JERYA�_�3�l`9��I�Q��eE�m�;ޮt�=+c��f�)��_�x^�R�Su�8nЋ�6p���Lz֊ȿ���򇚔`�#�j�¡{&��aR��ƔG�u^��_{؜���N�l�O�:J4��!��j�/m�)�B�fM������by� ؉0M	�m��5��J-�?�ֲV��#W±h���%�]Z3at�L#�z���a��/��u�U߳��v��(�G]F;�:=9=��n�E),3�E#܋���N��W̌�����5�^W[��úuL�M�rb�84�4L�Ґ�H\KT����DY��
�t�+#��~[�ukqL�d���x����Ǚ�;@��厘�`��V�
�2�	�<B�B��C���F����2�>̯/�*8�Vm�e�t_I��0��^ς���EM$�b�Uم��S\7q+h;wf����o<��������r`��y웊����o;ҳ���[�Fp�o��Ű�*�8�a��g]�!���a�� ������ƒ��)�1�,��r����-�A���\?����{�<�|�<���ٿѥ�]�8r�^���� �/�6���͍r;V<ׯ���'�l�	�|�� ��+�c���ؐ�zWF6�?/�	���{f�G1P0`���k
%�D+��j��xn�q5��CH�RtL����y�^9U���r��i̙�6K+[s�P�7�"�e�vA`�p�����K���Sg�J����!]h�%���N��하�ö�ve�19�E6��,����DTM$$ta����ә*q����mP�<�.;���a���d�B��ҫ�����꾚Cm+��F�u�
z3 D�i<-A���473���Hё�^�H+X~m���酢�����0e��ë��(��*��pJH�Z*"i�%gZ)ы>*�V�H2;o�֡PR��x ����HRJ(�;i�+�f��MI���^�#�p���;�ߑ��}���r`ɓD��;�=��I�^��]�[��X�"ď��z����c�\�Ǫjm+K��)ŋ_�<,/�N˫�.y��Q<�졮xڡ z<��#ĺYLO��`�U�ԜG��j���HS�&��I>�[|�̎qK��6��v�'���[ݰ�(����:�糈d��n����w���#qlh/ ���\W�K�`�`13.��,z<I:*�9�gΗ�D��	@��A摓l$���pw��Jb.�\�X�� G�bz9�ٜ���Td�	l��=�����X��ΚI�Ep=��Q������xF�n�%H�0(`�_��N�Ig���؄�������$W�>x�U��T��=1	lWx4�Ɔ�6)��� 濼U��������7��H<���%ny<Bn���jr�����}qt��]��&��I���Ԇ��kl�"*�/</Z�V*r�Ky�lU�z&�I*4i�캴O]�֨G��D�5�x���V�z�\�L���q��`�N�6<H$��g,���p@Һc�=��S�,e�c�D숸��x��\����	 ���'�������3�L֊�	�0Jd�Ş�iE�sW���k��Nƪ���p��5���TMm�h<�Q"�հRbM�W+Qu樂��A��;�!����j�ph�9D�r�X�����ַZ1 Q���2�o&冶ح���d8�"���K���nl�X-Z�������%��uB���m�M���z����-��p�x��Њu��nVF-/(Ym�������
�-��3���=�'� �`8d��`���d
���dLD\����Tte�_:�I��^����k�Eo��ك#��n����@�x��L���U����w)K���A/D5#�d���H���\_%M���_2��	vф����v�b��av�4�،��F��@	��F��ۦG�P�B;;{��ZD�t�z�����\��b�3�nHG9m��)}n�ً(�R�� m�X2����q�:�6��V��x�
h�^�=��
�/M|���).Ĺ�}�k�����{s�d0��G����������9J���o���C��U0�bI7��\��K�W`�u٧�u�j�m��#�Q]�sV��J�O�5;:��6��"u��eP����u<��1����ɀ����<FPx���T��{_�����;W��"O�[s-�12Oա@w_�^��#�;��)������q�x8��J�2�$3F���l���^�w�N�W&}_�
:y�R9�YV��$������k�[��w�gH�r�z{��Ԗ5��~�5���Ɏs�2�Q5s�I)h�(�l��*B�8˻�M��Z���kd0�C'G�@��u��CY`�]���c������eF�{X�]9k-����
�9�)_�n�� =t;�ѥb�D2�٩5;�L�0.G��9]/��D�� '~��x�)[�_�����A��T�h�3�tK1�������,/d������hgÌ������+�)&���"E����Y�8K��Q�Ȩ���В�����{�+|�fc�F�g���Bx)�=�H����{8J�* B��8�Iί�,K���׹�Y'뙁��w���Dą�8��s�
�`�f��H�G��Ub��	�ي�T@ �m��}�ª��4���e4o�:��4#�j���������ag���-�S$�Z�H�19oj���'�ց��N1�p�����Ik���D�%�0 Z���Y�C��#r��m�>���,C�*�n�$�����R
��Q�����{c�~FM����|�ۄ::��0dN�xQ��n9��+�xvv�M�ꎩ�w�Up�o���.���s.܆��u s�8
m��5�ƴ�jk��g���փY!�i!i��{r[w�,�O��'�Ac.-���P_B��,��3�8,�WV��Re!���t��t���͡��uQ������?ݯ��H�Lfh��%�����Z2HvI5�����~�q�S]"�:ѭ��� ���<��P�)�Am���������Pd�W����MЗ(�q�Lf�4eR5#�
:�R�)����|�e��=����t��E7��ԵO4�6�u2�ŀ�d,���p�v����x��.���Z�/��>�6H���U��2�&+1�&v�Q`���P1?������c��w�$5�l�୛�?�j��6%���m���s3#m��4��� �S��՝�����������s�>U/b���Z�.y̦�Wn����#�6s�9��8��x)*����(�J)�����(�c_���Fs�&�KZ^�T�j��)@�c'�-��Ku-����hL�0$&@���:2|���<�1u nm�w~�z[�8H�T�t8f.{�+te�²>��(�u%��p&���@/ܭ �� Э�ٿQ����܄/�ö��h9�$F��>̚>�1�)�WPqiM{�d*��4��)�0>��XQ*�m�#�5`��w5�|p�4�BJ�=�4�wA*ЇT�wĜhuK,XeSe��~��*�I���Xc�aѭȽ���hS�k��۵`k|������� �rY�-�E+2�نoj<T5<��Y�d�_ZFo�4����^3����]h���b�G������,��D�����A��fB������6<�4�ǗZtPV�����m�(��͂��O��V���(ɽ�n��qԵ�lG�]�+:�"c�HV�lEGp'�I �����)*�s���$�S1�g�f�M?5u���f���ݻ��S�P�㓵�$�(W(sX���?,�7�}Y�ܭ�}����<,��[��k�E�R{:ڞ���%�z�t�lŝ�СK�z�46��Ms�+O*���#��xt�[I��Ԍ��$�U 1u�Z��
��k�A�w^���c��'>��&C09n��p�W�����Ss^�f5~���f3�'����>@{��=;���X����LK/Fa��g�?�6s��|��+��aƬ�}� r�Rt�^�M܌�h�Gk)d" ��_��[G���#�J6K� �j�C�xTj����8��2�l�>�!m�5f1(�f������դ�A�������Z ��h]4G7B1[�d�8��|	���:`�b$�KE����n�@���ZUA\jR�"��D�7�_�����~W*)����*?�V"D���ey���{/�~L^Z�T��w�w0�	C�z�:���5�GхxOb����_�?QD���īԤN��Wk���q�X�d�X$T
�UC��d#�]��p)�I|��(r�F��ƴ��lbS���*UW�x��Xj�η}�/��(��ѷ�=9Y� }n�x�^>���W�����(���\Ja����Xb0�#@/3�sT�
��آ�]ҎGi�2�� ŗõ1x�)�uq@^+�(�h��[�+OI�+�|e�@�6J���W��W(�Q���M)�b�Җ'����p(�V{�7���>�ʽ�͸C(��4�$(��1L���kn��j�_lc����Lȏ���zZ/��(s*1��y�(w2Z��p��ߒ
/��1����&g�ۨ~�{ �z�m��U'_]5'Rᩖ�p�s���K[I�����i�=�2�2l��]�Gզހ�'�|G�<'�,�׸��\kS��8o�'2~a�pq�� h�gBKᴫut�.ȉu�y���RPN��ay��&0��p�X���-�����q�s������fE\�3<Ԝ��->��
4���$�������l�e����6�&�09,�7w�t�q8�Zb��B�C��A��X�ފ��N�.�1�r���S�GU7䤔��^��8���q�[Rw{n�s�!I�8��4��.|�A�үr{j�v<�"?T�HxE`����]&���S*�R�e ��&��Ϯq��E��0˵�t`[�W1U��Hm�{��ۂ������'���stǘ�mY���,���(�y_>}�'�2Q�5(*���g&�&N��t���D���ei�x��7h7�L��^����.�&@/�2����j�q��46N�2�f������Zk�qOhֺ|!��Ǝn��p&�z,L}r�>���2�6O�r�N�y!h�/�u��O}%^\�P��>%�6�CJCp�Cİ�V�J���*cď#N	�؞o �	�z��[�=jS^�1��W����g+��P��cŏ�Erp���scp�Xw��b���UO��Q#�N�M&E^���l����-=w�>N��!ۃ���b���h�y��=��\�7��>ҜL��HrY5b�of�n�k̓x�t��F�O���g�|�
���9���I[�_��y�
ܯ l֠�6va'ʰ��n��x�����2���qCyg]���v_p�wS��#6T���9;�ux�~��_���3�.x��d�+"ւ����-H�UQ.&��y~��@y�WB\�� J�;��G'�̜��&; =v���>�v3.��F���8ߎekB&�B�m҂p��~��}Lߵݲ�YtE�� &oH��9����N�Ɔ�����=��p�'~.�(�u�".�t�7�qL��	�
���*��l��?�#8P�����<��||Rl�\��7X�ʻdP�祢W������/�-�j�/�b����f�AaI]���n"'����ͦJC����J�3�����*�%0�Ա�W����������輵�s�b�'ߝ�)�%��B!��ӯ2��EX\ӣ��Zb�2�偌l�q"O{W�V>�P��h�J* �y�ݕ��P���gd�;�U��RU�[`s;��p��2S�ry%&Y�A�͚u�&[a�7m�g�͍&�o��D�rb9������G�]�l���0�"�[!���?ߢ�@j�"ʰ�6*4�(�Bz�Ep?��("$-<hZ�P�Е�*9�GҒ����#x����=*'�4� ��jd�m)4�a�ga�-��)�|$(Z�����J>#�y(�J7n��G�����m�aۆ�(�E��w������ޥS�U���J�<���(Uks��e'��X�r��B<E��G��4�o�v�|p�;e�U��4�Uq-�;'5�^�}��@Bu�+4�*(E�N�����H_����f���@���%�2�m\'N�_[b5aspȀ�L�D�%��N�������k����m��b�(aӝO%�'�R�u�њ�x�/�$�D�/%�<۾ep4X�7��ĈE�(��^K�!�����-w�M�I�w���w�n� U�,�3���F3��d���u�6�5��[��֮�X��"��)�c8�`���d*r~��tGN�����Z�6�(�Y
v�ƕ�i��ü�$Еc����ڎ�A���N��`RMw��ǀ�	m@8/rͭnQL�+�"�H�1sR�n�_���9��~)@�Υ]յ�n)[�c>#.���DrZ,�Q�9<4��8�s4-������'�hۊ���U܀8��\�L�IJ��ݵ�E�����D�E��?i�����	�1u�l��	xp�P�͓\6�4脶��s�_i)�f>�)���F��c�#���!]W=K�;,���=�V�\���Y�T���N�}i4�}�!)P�w�f#1t�m�a����ۧ͹�ܩ ]Yi4d��.��0��q}��M=�6|�,W!�DL�\�w\d���g>�]k�VP�R5��Xv��Q6�r���tK\��~�"��K��s~��h�],�	��9�o@�Xh��<��O�;����Gf�J��Vnd��Bg��MS�L�.�>$�A�G���(ӜI�5���$Y�^��`�=���|�W��1��������q!]T�$]���v�E>�*����-j��a��<?D:v@7:+�/�nL���D��f�,W�o������g����4�
'ɻ�L)�
��7��}�^��S#la'hA0� U������ֱ�Z�?^g�����u(UH��(�
]�^N
�X�OyVެV�q>�"��w��e�.O���6�z7mDߞdN2r�hRPy	B�x��E��b���["r�$�̍x�"Qϝ���0�aݲ9��v�V������{��l���RL��DƔk��2��=U���;��eq1�
��;���)�D�u�Ý�g���4�� U�V���%S��t|礥��P^�0��8�&lNQ�~Lhzb_>��mf˾�H�}����}��Y�_D�P ���\͜��J����!~��o�}��\���vС!���כbK8�gd���m��	�վ�^�� �s4E��l����+ĵ���>m��9���hF4u�z~!����=92}��Ӗ%)G^`����[dg�NPB/�%�T
�X��
�qF� U�+~ᳰ��S!�K�c!c���}�����Pc�0cl���L*QCs�����c�,��4�R����o��W��s�q+s�Ot�P�Z�v�� |��Cnb1���?���l�N$s�� ��h�2v����q�}��
)��j	a��s�=����D�2�V�+P�BKlr�qz��FA~ӽ/8�cNA\�,zL�z�Q�^��=�4���z-�����,�Zwl��ݰ��[W��ڨ�(Q��Ӑ0�*Uu("�K���W_lM�na� GPr4����}<��=�^�e&��(�d�������7F�a�.Q�?����Q�_p�#��!�BP@����e�\�m���hRU���7����T�!9Y���i��Y�glu�!����Xټɢҧ�9�ۚ��L8p�A�\�0T��N��v���*�ס�&����o7S�
�䌝�Z:ی�&|e0���]��fg�F���Y@I�7�b�J/�x�+t���m6�c��#T';�~��tڱ�Y�icem��������d3�(-�%�Ґ��5���$o�yYc���r3	��ʶ��{�\�{xL�s�����g} �~�͎U*!�d�hu��YP~��0�_
O�7w{��ʺq9L��ӒI�A��K͆�7����35>��W�*ݮP&���q��Ir��:�fq޽�����]
����� ��D�3:�G���97�5�a~Xi?E�5�����J�n��^;�ӣg����o�y�/?���V-����)���)��ʆ�U����_5:y���0��=�9j�Q�d�d�Q������ Օ	+9�	EJ1"_Sv[-�A�*�}i��97V�M�>kj��Wfރˉ���;�&�̓�38��ܚ�ֻa�\�j�@I�I�����MZv�t�B�Χ���9���/�����mp(�cq�V��������z�B=<���glGcǩս�A��0�V�l8^�ۥ����l+A����U�x�s��E\d�F�Op�`3��#a��b�?(����jtg.u�E쵮m�.����!?��Ā��;�k>��o�ެ���&Bǯۆ	��yE��Y�2�x ��3�5ܞ�plb�3�����zi�������f9�*o��v�����o��I��U�8��kYB���9�LC����y����2V��ʓ �9�^�Ă$M�0�vK���:a��̷>��*�RM�Z�i?��Ǟ �i7�z`����w���=ݮi>����͑/f�y����3��F���� �����p%���i}����X�ϾԨ)���v�O\��v3Dzt}���b��Kaj���� ��l�&i�~�`h��:o�	��M8w���٦�A�f8�H��NIƕLjy��_`H�#"Yp��l�L4�S)5�ti�����v*�}��AŢ(ZR�x��%VXO}�0�#,es�}sw��-K��q]�;J�fb��V������脥�=g�a��O�=[�&�U���Z�?�%:�#)�&�'=YDB����E�.�9_ <#����w�'�e�2�: �ī\�B �p7�����e9�pv���2�K���5N����f��;�=7�Yz#��z���qo}��M�i�枉�O˾jI��T��}�,1�S�^���e�k<d�1O[��ё8�D��E���4��R^��D�D?M��W&�d��* X]����4�R5�C��Xt�(���'!}������ K]y����6�ё-�@ �HuK�U	��'q�RoRmp��)��I�E�08�V�+ܡ��6E��PF���X7�*}s1�(�U=�|���Y�l�^�]M�����K�~���j�%�����"�g������pS����~d�"��P|'� �a��Bi�B���c�uv#�3�O���!�;�r��/�l�3e��Y �|p��8��FI�O$V�Qn.����dG��e&TVe�W�$��̉D����6�L�A���1��B�8��4=xp���2K+�QP��7@�D�/g"����.�ua=b��K�s�^��O9�� pQ�X'�aw"f?Qq`v���L��u9*���(�"�b^���Ғv�0� ���o���UoX��v"+E;�m&k�x�S�Ҡyyx&Fկ��u��g4��렸��Ts���"��tC-�%�ד�c�^�&o7��H 
�Vw�;��P(M��� u�:c��y�=0AVlA�&K�@ ���#�jq��fD���"���X1 �j�����;P�U"`�Nr�_Ə.)�X:�\M>o��g�X�����ap�	��6�mu�P�J�kk�С:;cJM�ƍ��E�����L�3Oʏ{Q���X��*�*�:��_�E���"�#�Q���kg���N�Le�`���c7v�z��>-��˟}h`�����-��um�Բx���T��c��p����%���w�w��mbK@+gi�K��6�zn��b(�����Tִ䇃4cc�_�M�n�&$+�`+Ch=�<�=Ck��=��ٖ -���_�6����/�NxN�]���!����J�B<�s��	ݦ�T'?�Q7go�ؓ
��^ ~ɂa$0u�enV��;��AM�rG� ����c��������s3��tUj3W�?�n�sS�؞<x�0+��X�\�� P:"($ء9��aGF�^�g�˻��ZSɒ5n��=�E$2P��,RbH%X��y|[�{�Sy(��q(��ҋ��¸ЅRR�L�,G��?Vj���� ������L�©���4N:�:��XR�����l}��`N�z�1����m�PB�����g��9�}5�{M7M�=�p�r���R	[^�o��(�L`��� =�|h+�z�ZpR,�ˮ�حE���}���@|�͵�?4�����^�b�{R$����2|���y�xEjDV�mpf�D�Ȱ���V�����ZsI��mt��~�f&�8{b7�7�/N!7�\�7�=��1�:1��Z��dW�w��T@���n�Oԁ���+�M�ڲ*{�0F-�D��i����X����W�������tӼ;���̓���W���e	K˶������F?����T�PמS��<�Fp�=�g���X���CI:�$\]����׽w��5���qV�Ml�Ǻ3�TE9 	2 I�����1��2��Q���v��k��)�S^���P7�<�!�U�[p��Ȍ��<z�u�|�3�߭���� ��V�zu��"��GS�2�cgA�����t�V��8��6$�s�h���^8Ü�DS�K%6@#x��uH`����ݽ�_�we��4
�<s~B[%�W'S<o	ަ�.F��O���x�r�SY26�z��>5�,<���� F!�W��܏N7)�8(���r~�*G%���=*A
���0�6+`z�0�˺� �����n�ZiI��3��ff{C��(����d}�6 ��W������"���j���T�hq�3%�s���qon!��6���Ήpl�,�[��]BCq:�'�x5���%���[&�o�l�F�GGƞ�=>��q�Xm�r�O�)��Y�O�kK���+Ҙ�*�<��M�PR��ި���/P���g�ۏj��痢�ѐ��Dʨ0���g&�	�烚Ne7AyU�x�E��x���ǹ J�
�ݙ
���WB���D5@��1�c�na�*(��S�2��i�<0_�m��Ԕ��#]��Ї]o�c�O#|0F��s�wq�"�a��x��
��7�IKũ��]_�H��dO��?0�q�M���M�*����^�Ra�'�0�!�8���2�_#��\�����i1y��
�������Wӛ] k��~��NL�<%��iѪ�x�����B?�.�%8�8M����t2�RU�5�A�'x�>ӟ��6+�O���m-��i��%� �	��ܧ���\[�����刪`�A �Z��:��Ҕ8���	�EΈC�b:34E�� a
_;I�W�,�e�O���˵��Q��xD�I�&�$�I��Gj.H��g���8�s��ua�����F�2l���i�p��m?^?�{��E��{�Β��Y�1�O�,���� �q,>jg@5���X�сGlH��k"�򳀨#k��<�^����>RJ'��n�P�+���'I|�u{�f�>K=��`M�� ���W��@8 ����^I��i��B�g��2���sPk?�&f�� �������#�r`��>��uywrE�ێ�d�q��"gV��lM��}q@��C"���MT��6s��X雊Σ��]ĸ�X
�KӺ`��`�9�3��$��ў'Or���ǜ�*�gَ�	��d_y~G틧� ��-稗�vu�����B�
��-~g�d�_a�%!.�	�K�Q��
��ZS�x6���<bꔜ9��� ��4�@�������W����Ӓc]V?pe�=��m�p�g=a�� ��y�fS\����M �*��8��򐍮�����+6�)"d�����M���ie����h�?ʹ��g����Q����*��2hXx��H�+����+#z���4!O���5��H�[nv�fp�9a�zz�� z��fXc�誦�4Aғ�G�N��?�O[��*o�c�Y:��q����`�[d'A�r5�o�|%���������$��L�����O<��Bd��8!֟���-hnE�Vτ�T`�Y�y3h����<��BN-�i�,��+�h^���j�k\�X�X�Sg���]��?�31�w�Kcn�[�1[�G]�m ���}�����4�i��B}o�wecd+QB���q���d5H���N�5F�֘=�I����<�z!a�֭̈�:��a��P	����I�(�ug���c=N(�ʱ[����I��AsI�Ǒ5�3� 7C��_Z0��D�˴r�M���\���)����{0\10����[�ȴ�z��m�d�����B!�4�(���7�u�FWc'�� �ϳ;��A��mPW������:C����� j���8�t�Cj �%����%o~kZ*���h��ۆI҉.��.Z'�2ܿ�� u�سd�Z���8����$��[~�]g���g�KC���r^sl��¡����V�+;����N�.40AB��7%�u�2G���������¸U�(��}�̉L=\��X=����(%�+VJ����L�/��#��Ymd*�'2���	�o'����&��nC.�+N@��oQ;>1V:�Rd���Ėk=���7~ݚ�lֽ=W����!eW.�3���%P+�ܭc Vmm�k7��8U<�%w�4�M6o�Z��/�y���L<�|�dO,�zdp>�������dUū��4`d�/�'Bq�Jk������!`���o���suȗaP.�s>��pq#�1��Qɋl�Ҳd�x
\���E�e�0Gakĩ�j��p5Gs}%���͘B��Xn�m<�d%8�,�>Wd��\�-�q�߿�j����eī�f�B�Za�t[��q64���ZӒ��\[}e�`�F �d�a��R����o����cN�Rd�RJgZCb��c_�:魬f?�3��Z���y���8J���}����A���C�Sm��w^#����O},}�b"c��B�9�K�jÝ��6@n�$��
,X`���֠�󳑧,��W��m$
�6J"������ox���\ҍ/��܏����:�95Q�	'֬�_��+VX��\��F� �W�/H���T��;��aFd�)�����e"�ܷ��	�z@j'Y�K	V!���8�;~`����
�M�7@k��C���a��[�2}����=�ReYްu9ؖ����sKNr�p���$;<]͙�%~A�U����b��bsv)�7�]s4��f��Zc�v�������	�aBq����f;�Q'�W
Љ�00�!<6�zD�_��Q�VC�����!y71ɟ{����2a�ͬ!ǧŀ�����o�kL����k�����#�Ԙd�4�������؈�k�c{Y�7�K��@��XH�83��@�Y�*�l��-�����_����>�Ȧ�nVteѦs��*D��I4maw%�F�p:��ld5�!��˗t}c�vVj~s�/���V�$ɨ^/\$=	��5�k��NX�[BKk�0�@F�M���មRܧ���Pک���*,`Y�WJ��ǿSU��<?Zy��!�a]{- �qDʕ�Hl��7OE���z�[f1�1����$A�}��I&��2�WS7�*0��Ȅ��It��qb�t�Mx!-��:J4M��r_�D�K �>���ٗKy�<���q4���F<0�©	��J��Og�\��qr�#��_�&��q�����b�L�|Ԃ!�)8�`�>�����6XE�m3P�}T���ɿ������_35�rpH��S�aHg&x��`Lw�5<�_C�ۚQK�Jq��o�M�q��̝�N�$�>&
a��<�::O���b跊�������zKl 4�̽�0��B������r7�6:���6d������x�	=Y��
��v���9�To@9iJI�a}\�H2�ޱg���T>uYVUʍ^Us�Kpy���{�o�&�P��L;1n�B}�-�,2��H�m���{�S�<�m�&����|/������$��֭�	y1�~�+g�_ipݗ�"�z��v#\��+n�b0���/������#S�U^O�^��x�[2�����dޥ_��SP��GX�Ww0P�͑��:w;��(�Ѧ A�#Yb�B�����L�8����q�h��{�8?�=�ӓ�,F`KrL�O���h}b#jgD�yM�sKm�@N����� �H �� 4�Zi<��LRu�=����L��T�f�i���i=nX��Vh�T���;�yph*��eHVlԈ�(1P��y;yj�?���!;����&~k�xy��ρ�]��HQ�N`�_���A�l�ҕP0��f����"�%NS^rR��쨫�'2[�B*��[_$ѳxhpnE9k��M�n�K������/GJ�ŃT\̈�d?W�9g�T{N;y>W�( �ϓ�RK&d�vn��D����BV7��$}�R䖇Mn��6���\$:�ń���
uY/��V�'iíKx ��"��Eu˅k~�t,J�b�{���)���p̯Pڋ�
������2��n{o���1�6��7 5��mX�d�����n(f��d���
�,;|s$��/��`"e�pu��am�	H�ěށ�(޶�Ǐa~v�~��.��u<�Vk��1a��0�x�p�'ȋ�}��64\�>뜩��ޣ�ϳ�%�sK�˴���X�0&�_�}Q=R���"1n�L��+n�n=xpv��%�k%���j�5��#��-%��e�٭Lc�G��������*~|�˟K.H�"�l��O�_ny�����T�32f����c�,P2�=v_vb�=�8��C��L����&��0.4+���N�_�Z�Gb�M
?�ֶ~<�}\��^�V�f?��P��� ��.p��R�G�Ol�H	���<� J�SvpZ�Y*TP���Aew�p����`n�n9.��5���=4������9�Yá�S���ɻ�T��"�_����f��yvB_�Se�D�J槌t=���l�]�t���C0�2%6���½��e���\�IOMF�$nZ��̥KEd\|ٕVĚ1@ו��ee�Y���o|ʌ�sj�X���Ff�xM^���b엪�?4,��8>�N����N�ĥK�vy��ϧ�eK�@���~8x���h���6q�D���Xc%���__y���<$)�Ѷ���_��.�9(�ަ����_@�!c=B$&���y^�T�?
Yߓ$sĉIH���h��������Z�g[�3�lo��\K��\�a~H	���?�թ6�'�����5�9+\c��k�<M7�
w#Yw�KG���Xfb�$a��. �3�@���C$��/�R����REJ�Ωq����Kki�~�D.����%KP�
�;Xo��F2����h�u��t���h��/���jG�<�iʧ�����Yo�G�Eό^���*W[4�@�ܭ9Yq]��*�>��5e�Z� ���DSf���}�>]�Mmr���C}�~�F���i�=QLW,i�J�BGw�2$�ۺ(�{���b����<)��16�\M!��G�1,�\*]�M�L��ʘ2� s��$��_�$:�}��G����[0��6�N]�ߣ�S��f������@�)��*��/u�6��
Hi�(���M� ��i��b)j8�����U��cLU-�\<���u'�����A�192�����8W_ԫ^��XX��(5w~��׀Nop�#�����gJ���^҆�WK�r�1'��Ӌ*[#T�j�Ӹv�t��߀i~g��F�8��:�aM�D�����lj���#����@j�`ѣ�c������o�Űm����f�������GR3z��/�s��b
{rU��b���q��*^����gح�(���qi�jN_�rˍ�(R�Q��wf������.I6�\-iRcJM7}Z�ba�4�c�Q�8b�2%�G$e����=�~v]��Z
��77�z���ՔJ�|��e��[��N��W�0�4�Α��6���/�*\�؆��x�H�f����Z��>ʶ����_��F�d�jF�aߔ�Cd�g���=����7�� L��c��?J�6ƍ���1�	�S�S��`��ȷ�p�ť2�Im�)��U��3Ƶ_R����\��s�w��j�Dw<}�C�e�Gtſ̮�8���5� �tt�Rwҧ>���
%t;f��ȧj���"$ս��˝�������5�N<�1(��o7&�w��$���<9;�HF�4�"����l�P�Ip雴�V�6��_Q�-�B	 ���FS��Kh��2i�(������Y��g�z�6Sm�$q
[�J�򂗅D-�5aD���)����#�\��m>[h�C��׷�\���R=���/R� t����O���0��T>o/�o��(Y?�L��`��Dw�d��k}^�E�\��v2��.dwOA���f���q��ћ
�84/���s��3ASJ[��z]m����ڀ4l���
hO��z����#G�G2Ȏ%!�8#AaBM�z�W�e3S��%�B�D4b!�0�%A/j>��u���bI&e����r;�������?����G��]JĿ�z�C~�~9�
��oK�IhP�ؐG�����6�)�{�\������W��@�����St�J��pZ؄��X$��?��ҭ}țT!t2_���}�ܞC�2���f ;г�Ú2S�2�^�Qc X'�X/�2�9�'��M}l��<��*�=��H�Bd�G�0wb��+�M��{1���
bvA&*�`��^ύ��z�@�G"p_�E�"6�KH��U�4x�I���Ֆ�������"���	�B��Dd1��$��ƟBTO��$�b�Un��kW�+^��|^�xu��P&�yK�{�.�w�D��h[{7��P�[þ��fQ<��̎�Ăc>7��*v�.�CI�{$�\cT�?�de��� 0D��-|�i�D�_ 4�R=�@�?�žn�?�O�V�4��j�{m��l5�0�&RW����p ��멾��wA���r-���v�䏦����Cl̓�И%z}U3�$x�v��Ci���:�mm��]����լ�L��$�Ԗb�����*��W�C�kD��	X��Ǌ�4��kz��p�M����r�㶖��"��QF��NMB0.�3�]��_�x���Ϭ���Bd[v~'[���01�5P��Vɢ1�.�����n�yŔ����^���B�3Q�&���B��&�j��&Ș��1��+T�y��c�0�1��kA�Ѹ>�''%���,��å�ڦ��!������~��!%"��g�JCk:�����.� 5��>9Uh.Mx��Cc�Y���2#���X-s(�O�E�	!DX���HW�Ԥ��P(����_9$��י)�;�1�����X��{]�\@���0�2ʼՃ�&�«�V�^��'�Z�ݎkn��t�&�?v�<d,ωGh)A�$�{υ�ɵ�S��_�#HITU(�O�
m+�v���M��� ��|l2����f�N̏�Rp�dx\0�|7���A�xcbp�w�ۭR3Ǵ=YP�5RZޱ]<-vqLˈ���]��B���]6�%�m6�)_!�_��_Y)��_���"���z_��5�㝶�$N^��`����i�����ԟ�
&E�>��)�aSNF�8�ǞY&��)�t����l��pKqz�\���ƙ�r+I���dѣ��l!?�Tb8�y�/�ĿԘ��Y�&�� ��L��@?_��4��X/� ��#l\O8`����44�7��.���P>���c�?�ށ�bi�����%f����(����W�)����ϯ�&C�:E��`Dk,"J���_�a������5�e�}������bC�!L0`�X�m����j�Ak�n�v[�����ԏԠ�=�NMvJg�u$?S���~�2��)�:��0:P��IB���z�̏�Q����ӂ]o@HKOk,?BS�:	�Qԡ����G0�#����Ȭ	@���9B�K�~�̱�r���Q!���<����z}�H�Hg�����6�P��\Bɽ�Th�b�.�%�����P�U�Nu��:����:�ZJ�vf6�o�1��� 8I�'C�d��k=�a�Ԏ+M����>������'д�)�~D�/�M��L����"�l����AKӨ��>�9{1X���7�L%�3�\�e�VL%��*@}���_W*���P��GZ^񆂽�
��2H���/�2��H=,�������+��h/ŰsP�d9	�!S�<��sH�[|�%O���ڤ��|�I^4ea��@���1R�=AHF_�i[�g�&`H#�繁�V�1�a�{��x�Fi�DL�rr���h�I1���-�˼U�P��t�%�j%o���4ĶҔ�~L2U_]%��|]��~�0¦J�I)�Cb㩥�ik��r&i���)ʹ���~���� �v�H�����>�����f�S	�i�`	h�]�_T��p�/�m>�E�xWCP5&p�_,*oJ;��^a3"�z�	*f̲�ݳ�Yѩ狗rӉ/��;��6e|�v;پ���W��?c�Ƀ�Ls#竩<e��+>�<P��'i�^�)�y�~�|�]���S�#U��v�E.UVӔ�n{"�丱�ɘG��zE��O:ee����x��i��a�f;na-+���?��Vs)���-���gk@g�_tޅ��a��`L������0��6�K�Ǔ2m�:ke�@��#�!�V�w����ܸ,���<Em���Jh&��Y(%$�t�+w>�X,M6i/��)6_B�̩�}�sR�+@��l\6�è����2�O�gD��lQ���v��8~��e�Z�&�#U/�\����	3�����46�i�vm�߯�8e-2��HbV�]q����K�v+l��%���u�Ge��~�.=��G���?�����<,�����5�����I2��U#��&CK�В���'L�������EIc��m"u�x���G�575�j&K�J|�[�#B�-���P�3�9� W���b` ����GTOY�X��V�K ]b���x��*�8�v�$S �N[�����Ɵ4�B�n-�t ��<k��7��4e���n���B�8�c4LgS���� XVI;1��.63�#)��y�Ռ���d|��.�����-����U��>�z����@������]7i��������b碢ڷ�h�!�[`S ��dT�g��&OQ@�'�� ʛ��O�9���=�?v����Ap��٬��s+��@yp�n�����(력�=0�%�:h#�B�����^K�fs���i�"Sո�)b���{��C����v̿�Aͻ�c��S��?�F�Ȁ��rct�U�d��}p�5?ls9���į�:f��wa�K�	m	k-�^uB��[�ª���t����H+��Qz��3�3rʅ�'�XB��aK�y�&if@��u70��F��F��a���M��T��t�A���C�8�t"W��Ë�с��RhÓ�z�M�Fa�A��$������>���9�/K�"ۓ����h�Su���J�]^�c�'�]�)ݐ��\�l�n�M� b�qH������e�E��Q�P��c����v�𥤉�V9�GS���9OR����4s&,Eܬ��﵌� ӫ�u�&{�^K2im��>��F��m9�@_g��ɦc�����VX�N?r�b�M���͚.´S9QT\d:�6E"Y1���#p�����"�9��zN��<�Sz2�ǔ���@ɪ��c>� ��3݌�S��%CE���="ױ,��ي=�����mc���h���4I�j��\��E��RC�L~�[X|���tۑF�i%�Dj�Mb6̏�R7�^s���XD��������g2_^0�Au�y���l�_]L�*B��V�-3C�Q�[��3���j�x;�b���f�w)uSd������gG�=�"}+u(��~���w;N@�Sw73��,YS?rCnT8�Wރ/oc,�^ �����jJ o�HO���d	�\VO5��92����ok-�� o;x��8��K�Id,[I�M�#���A���0(�t�gG/���}�=صX���5cy�x�o~;�n����x�wa�=��Cۧ��O-+i𾐟�%K�G�d�Mr2��u)�����NL�t:��S��cEoT����@�)X�+��������{]������<���9 ��gU�"�+$�<�.f�����	ys���gUKh��6���ҹJ�!�;Y�~-�Z�"��O�����!z8�&�s���@ÌJ��*d>�X���g��O-^w	c�U��%�+��tI��J��f�M��db�1	p�d�Y�s#�����.��d�:�#�.
�����7X�e��n�[H���+mU�Xz(�
jLxG��*��[m�MK;�����U���y�}7��z�?�U6g@"�7� �죆�|��G��i�%�T�Kc��ߌ�c�̱w�AHϧ�h!go?=~�@����ߒ�}_AA��[���<b��=�`�������:(Ku����3< ]��=�V�ls5�����+��9���#��lZX�����Z��D�20Ϝ��$'%��^�a�˓1�^��2'K�`�Vބt�?�Y ��h+�5�ŷ����FE�M��w�; ��:�E����һ��W�������PV���Gq���K�`�+}���Q��i)��6'���p��O�/OPw�>�V����bR��[w��(/��*��SN;wi
_�=QfJum#|�J��7��/Y�{)��[�f��������M _�ژ� }W�\v?�}���+q[��m��X��kN�M�T	��M��*�/��5�俬f���a��B��r��nmv6d)>S�Lx��	��}m�zedn}`V�������/w���
���Q��v54�[�A^�1!�짎�E�Q�>OD���P�}��g�>�P!�Y3V�E-ծ�ުK����tN�x���|;���xq����������=V�G!Q�y�x9�sK�6���B${>�E���5:n^ꑈ�fv�~���衎�@˰����O���#UD3���@/�Sc#d���ڕo�� !���`_�/K.���u�n�-����t���`SQITت�o���+cֈ��U1U/�;>K��x���D�?���	����n	����	S�������՞�=��P��`E,��iO\�R�{����B� L���΍�F�O{�_s֗;S}D4��9$6ӵ"�w���3��kK+�%M�|����cKKc��Hĩ����4��C���َ?����V$hڑ�.��y���t���*����A8"`�-�3��v��Om�r��ET�AR�A���0e�6� ��1Ȕ��N`���T���:+�-�F�� �B�A�<9ɼ�S�f�k7�'&��ҍ��F�f�E�7(zu[�o����$�����բ*��4��3��k�����<1�~4HC��1 [�H��h��1�ҺtN~��/�����8��3��&������G��4"r^T���f�s�pw��'�M==�~7�����M���=dښhԡ=��:��\$�����stL��+y�R��8�ɴ�ź�7X�m��/d$��+k2\�ҏʸ�	�m����$���Y��mӱL�iz�+i+:��j��y��1 ��?�e�oK?�5J��gn�	�ˡ��\9���>v5�����6����w�׋�͚s���5�7�`�LR��0�7r�|���t�È���W�IlaǍuM���)}y�����H:T_�?C�I��G�.�;8��I0<��ۨ�hv��4ݐ��{������5�_��S_6�(`�i�G�j�6�%���α�,;�w2q��	5���s�ቡ�'����bH2��/L���Z:(e|Wg��U��.3��~�����C^l�U!VUsS ��8}����A9=��,-W�c��fB�]�+���
t�㖊���E��s��L��=�@Ӂ�����et<N���dO�,X�$c-�)�8��`g�PS���8m�����6G�"�"pl���̴���׆J����ڛ��q�F!&L9�aٖkyΜZoG/�U�J�L�`B�v����Odri�W��{-�)�-�tg�2��o3�Zȯlo#4E;�=�/'_(Y�A�wy6���ZB�k��ɧG�<���1v�v^���1�X���
4q7Ĉ��q�uP=۰�Y�9xl:hE��~�`=��d5�>�����*P��
�L�)��U��JT[<�T�T�����HOOJʃdQrmBY�Cؙ�����^k����}�7����d0g��t�o�!��4�i��q����&�-{'���2P�K����Yo�Dv��~c�R#h����Łnf�B�7̨���-�L��D�F-~�6�tJ�4��y`6��,�$$V�O
���U?>���#�ʑ��})mWP!̕s�4`jG#��`���g��ف���oo�?���Y��^�f�h������x�V#;�);���~踿s�=¹��W�Y!¤p_H+�<�t�v2��>�F�0�ǭJ����sň`Քǉ���t~����a�6�G��������M���uB�⊫����@ә�FVfC�3±!�0v���M��:6��$&�D>�+���3�������{�4������up�RV��0�_V�F�5���Ki�!E�`E "�����'�A��?�M���YH��s�. ���Gk~
��H��eFo$׋�5:d�����9�s���t :�zv��Y�	hW�/��{b��NyHʔ �FM������hl�A�F)��o�ky98���8�z����u�Ȉ2��7c�n�6����e�Xb�<�x����p����Y�����{��rdL��oHq�FJQS���w�zbSp=O/Z�&�(y��;�<ANgTp�5G�-��x[u�������掐��յ �+i�7/W,�%�� A��{�ee��Z���7����z
��D�_a������[�	��!��%�Z兔`T��EC��o�.��jRt���}�n
I���[��cH�����M4�ݙ��p��=(�R�Yb��7S�� �k��j
ތ���Qg���b%t\�J�
|�*��R�'��\�J\�Ay�G|���|�0#�Eٗ���:�|����l
F��Gpj��rK�Ⴣ��@����|�C�kw�@���֌��_�ڳkā�d���r��yB�!�,`E '叓Ń=~�a��:����	�Qqi��lz������Ĥ!�����X�W�ս�՝�7�s�^o�`���*�����J�U�
�6����"�Z W�{V�+�>�����>B<ޔ�q��E~S�l��,	�t�`���c�ddF��Z"�6�KL#��uG8�&��+��Ѕ泗����A�;�p�eS��Pu~1
�i�1�(� x�%zKg�.��Z�y����M~��]�Oĥ��KeetN��/�i�!/)��0�,����,�ȋ���+�oSQ�f����%��j�����»�0���]$���� j^��~�E����[{�0�̫��\I�:��2%��"��D	Y�+�l�_�
���8!k�5�.#��h� d��p��i����#i�e�=0�c�� Mt����n��0�Eh]��Q��uE&�&�X��PU˗��2g��5�WC�D�׸�����1D���QۯPBhK@���˖g
���9ڃR>�v�8��.�{��:,J7BY��.����HZө���Y� ���$�i�_�@����E�.@��O&�Cna�=R��(�_{R��H蠟$︔K��_����m���W�(Fy�*?�8͆mfR-�����Y���f�Rj����S�(�Qp#�=�p��IGBx�)ظ�c����������VR ��0����^6���[qy��;�¼�v]�{��LNaǭ����<|}��	�(�������f�vo��.��i`��$�LXǥ�*}^k.-�Waӆ�iuzÂ�.e�UYB��a���?�z�.�A1�y�@�����8`��9c[�?a靽-N;�q�Bx&���G'T\)5���O[YW��U��0V�̓I���j�qu������E1k	�:M��v <I\)�U6ik�0]6�{#]�����{�ݿ'��[âYl��5-�
M��h�-w�ګ�'^��[h1)�%����) 	�}��׎&�x]�2��Y�	�r%�����u�����������3�@ӏv�:S��_'2�!�q�#;/��O�9����Wa��j��x{]/T���$ ]:b"+����a�������=$6� ��難�=�/��g��A��-�$�G���ȮQ9� ��\�������X��
�ZC�
��c`��JiM���K����#dS�h���t-뼃���U�&��2u��/�Y�z2��(�.�����4����k[(�#�E!'�:��G-:L���ws���'xJ|l Yfe�c�G�B�Bݪ8����z�s�AAf�c:�����	SwKٌ�R,}�/S$��6���5&Vq�Q���&�U�A��^��ϗ];�G�/�S��+<���ubI
�7���VS���>�������|��]
yN��bh*��0I�RŚ�@Y^-�HP��TR2Ⱦ�mZ�}sGZ����Gn����aQn�. I���)G����ք8�
����Hc��{��'�T�p�j>�ah�;�=�<�Um1���j�pq�̮������dA�M��I���ѭ�����J���%vjG�p������W���a`�9�&��a7V�#��O
t�GԎ��# VZh�%su�)j1=�m-���)u�hM���L(/�+C���p�~nkc��	jO���ۨ�v-߉�I~� *PҶ�FN�%�;S����`u�T�;B��h�M�)�O�*�{�4�=��!g�7�z�U��������<�=�_��t�����9]��2ΙW#c�*�78�733���!��M���cW��+�GK&�]OZC�<�z�OBNT��C;�M��;����6�� $!�gc����`���3��NHwp�q��%jR@W|l��o�N[hWQT���RY5�⼪|�H�X�r�����?f�<3�oڠ�>�7:�����,��Ċ
���o�����j��� ��^Ԃ5H��@����-	�S�5S���覣'sUn���7,s����}U��L��c��Ǽa}>O�\��`���;��:ø��)TȜF�w�ԕ��9Yp<���b��.~{��׻�	a�Wd����C�(��k�W�jNvOU�N�'U-TT��+�V�a"��p֠���f%����cC�k��h�^P�&��.�a�gd����v��8V���
�.0�q޿|�n���s��ԉօ�1���b߉�7����\`�,��?Q=N���Z�.P�M�*�̱j�J�ݜ�˰ %R�w=br�/��n=I>A �Fn����W���Uj-�ƶ��K)y�,�o����,+ѰhL	t똟�����(�U$:S3kdb��aEk2	W%�D
M��������~�O�C��g��o��j�eP�>Q�O�N�E�
uit]|��$�w�����b���9�=�`]���1��5}���jQ��\e`������B�+��LP�6�Ɨ�3S�uz=���ֹ�n�FF���J'��b�%�;+�!�tj�n�TK&�(�'u�y����mw���~
��(7���\��d/h�n>k�«�+"�������J.K|+O#�����#h:���xw;�.5]ZwIZ��/cn+w�Z������9ċ'��F�7�P(YN�ט��O�mb�w�Ѥ~��ɪ|үQ�N*��O_P�)N{y�2����sH�|#*����_��	�D����˦��W�U�� ܆7��QhW�� \)}�5;bz���)��	�k�w�hc�*�&?*�	7y�?��4��p���(I�B�+�˵�Qm@AY,��9+ǖa �59ʓDZ����;hԛPJ��E��k뷡��%/���v�k5��y�L.v����u:w%.��-���7�Yn���|������ݭ	(����m_���܋GఉX����a�#��jnɆ�UŃ�C���߀�z�"|���K	���s�g�fU/z��ł��*C��^h+5\!;� 'ɍڜ)�x�m,�K���z�W"1 ߬<|��qy�;	���tZ�U�heZA�B�_��k,�==)���;0�8:��L�|@��8�wuȸ$9��P�.Cky8i��B�z�ˇ���2졞��k�?p���r�yp��{cX�b��pB�{��-L�A�K��7�R,��	�n�R��'1Ι{Pg㊦��AW ��:�*�5�ŽЋ|oV����~v7`��:��﷥�Tg���1pP��SE{*�MJv�p?�h�B��n�,A�k��m��U%�?���b�!j�3K�9���3Z���3��ok5������"�.����N�fJ�ׁ3.��g�$���&7Fk��^�劋ZW�,�MbM�Ĺ	��Clo�?譠tw�2"C��%�����BЁp� ��<�"��.����	���MK� ;bE����j�j��k��t��g���}�u�C�$hp��RN�lI��KK���D )wd�43�H�3��|%ͤpx�V" �_�tIs���
[�ڌ�u��:��l�t���.ӰZAu���� s���;�OǦ�y�%u��lh��#���#�W��ǯ
p4
��Y��q��Ed�/d<y���th��y��-	�K���)FX�\5wb,}2-ˢ'^WZ!���w��D��*��P�G�a��񅝻/�6C*ݏQG��o*]N��m�C^�����Y
^�S���
E��z�{sF�RW��%������/��[A�=6�� ;��}�\d~5�،�[��-���8%"�p��9C���6��4��(l�Fr�B�"�����&[�j-�0�&�E��y�u�*Mfq';��M�a�z{T�A��ci��/0f���g/�p_s��"m;��gO,y���cbM���2�8|܈�.p���/��=�lu2۲���ۉ��7?�jx��?�@��Y����������z��˳	��d��,>�G�[oCAo\XDXB��Ķ�,p��a�k�m.!�B�t�ƎE��2�T�A�����:啠��O�Tz<�O�]�Or�uE"�G���Q������#((��� U,����	H��K����v�����hi�5�hMȊ�#v����7	���$�m������ru:m�<�b�~U�f�	>��R';ֈ��h-Y;xF��v^�d�n�Z��oz:U���L}!3��T�A�X6.��σ�#�F�,y�-y�B�ʬ�[4�j9{�7t�B�R>{O�������l�����"�S�^!��R%p���'�!W�CB#���<q@�;� ��J;V�����? �mH�q��2���&+	�S��j�;hɥ��*]V���s�k�V�0���gӨ���F5�F|�Y���$�%zb��PDt�4��5Ag�h��Vp�����4#?)N���Մ�$��p�~��5#��7�$�-��k�@��^.���Nxhd>�����	������� ��ӼU����X@��k8���F�!�s��7OǦǸ)�:v>D��Oq���qDsj��)ihmȚ8��t@ٿ)���&�l��@$d3�̿�޿(���Wr�˱~��*�? F�n~` y9���2�~�������NءB����c_D�ҏ% p�\6Ѷ�w�tJ݄i��A`�Z�9�}�m�GC1��j�a8(�v�?���ڛ	�k��o,��u��ވIG��>����%"3�[�����_��[�sA��ujn�XP�O�n�XK��j���x^�(P���peW����30����2�q�+$S�"�d����Æ(��u�@��7}i�C]����j�\�����<3���ϯ�P�ǻdP��X��m�Ä�M�NheH9�Dx��?w�+?��ѱ!պ�
�R/>}���UӐ�tm�۫'��G��lO�<�j�F�M����0��MZ:��Ԗ����Z�pL�M���l��k���t[���3r�"�r���=�;9��k!�u7�|^J`}!�ͥLB������Bw\B��{fe������i���b>��3��i���~L6.I8n��c� %$2�l�w/�9�W1��U��Û�Q���x���^K�BU\L �k�W=%T)�V>��_%�S]���^?��O���6��!�kac�*����d���\	���q
�/�������8qz�'4�Ǐh�*O�taj��1��6���Z��f�f͊S����l����My�0%t<;��vG��}�"����� Y�]��iೋuuqN.!gN���>�~�RXDv��v��:��ɠ��^U�u�l�z)MOxQ���`�����BꂄCE!���1��QB���2ۍf��:+���o��i���GX6袾K[���О�f��OeA:����ԛo�b�ޤ�V{�~0VO����>��;;�-�-ߩ��B��R�c0n��j�"�9nE0�eǧ/��l�A�G3MǕ}���y����yJmyaA����iOk4�RԖ�8P���X|G���u*�
�O��ٍ���ͧc?B����q-nE^b���-J��5i>�ԑ��PG��Ĳ_EEVyŮ�,�����زL �t`�%b�ׄh)�O�~�Χ����rሀ<�6�N�[XU� F�P�Rr���,T~vX۲ da�SQν���wխ����#@��WD�`�o��?Ud�gP�KfE��+���e[��!׽��m
8)(�]
 ����c��m�c37�?���bެ(
,b��4��$v'H^n0��o� 7�M�X(w-$9r|p@�G����{�˭yW��s�0��)�c�q��p%R��j--k3���Bkv��ê�B�YT���G�Y�YKo'^?�T���v�> ��ؿ�w8�K�����`|hO,c���*���mV�t����I�D}<��r Ny��W���_�ƽ�9��-����ٲ���V7�:�:�ZH�Ԛ	��K�_�uW���K=K��%��*�ᓪ��C��+?-��T���	v��n���=��90��P��f��2K���x�-�����y��aȲ��ǧ�h_YG��׸���Ky~5���G�6Qe;xjh��#ڗM���8��.��E��${���@B�3}�T~N�)����|�;�N���iʲ|�4���G棇&�b�S(�ɳr"7���`��,�I�? ��hPIc0�D�Gpnv�P���c�!Ғ^�7R߯�!��&V��_�P�v�ß��f�w��iёB�V����|p�Ӥ���Y��s�	���4�!�L �U"u�'�T����|�)M�hh��ї�P�cK�m���r!�F���
�����	�<��~+�����
��H5�Ht���geXBٲ���]f��[Y(U$d��s#Qm4�ܳ�F	Wv65��mM� �# ;��3��"
>@I��
�P"mG�;&{?Lu���L���=�8F�T����{5dMD��F��|:��,�}���1օ�v���K�A����t�^yN�1
�!?��/�r@���D�K���4�����hv��b�\���,���@g"`���l���Cf.��:~�"����r@�����k���AY_#��~�G�A>p!��@oEx��;\(��9'^K���:|^K�!~
�sd�����Q�}�������)���iܨ�	�,�ؿ=ܮ��	����7�?��#�6k���J��������wQ��W��,cś�[������u�o ��L2�
H���� �-A�|�nR	�-�\�r*���l6 ���6���k7|����g��K�[��M*^�$k4tTD�y�8S���?��b��⒰���Wr3����뗳�}����{�f�Y���?R �߭\��Cϲ�ˁެ�P�O�O��D�Xf�^_��C&�y���9�dh��Fr��#�Y��J��F��R�X,����0�.�s�έ(�x��c	w"��j���y����Tc�w�-�T�Fr9��y@��0�,���h��V�m�]�Lmv��\��?�-?:��̬�ų̴�)�#��f(�"*'����9}���a�fI������Qp� tR�v&��B�b
L�n�a��gʦM�Tł�'�n�t�FC�\��
L
�0;�o���B�3�m�S?�x�!|�V.�\��S6��,�� �^�����F>����m���Ԙ�
���@Fr#@����$f��>f|@ݽ��*_�_�1��F���"�Gg�Cy�������1?��<�?�X�D�V����#$�Lu��N��L���ᅎy{��KOq�-��~x���%��>ğ|�'�$c�`H�Y��TX-Ev4�lR����H�����dp�T��2�
����"�蟒��d)^(]z� ��cF1��Ǻ ����`O�J��j�[�*��^�9���hd����ߴ1qI�|��t '�%v�� o�t�
�+f,5g^���Ds��p���݅�p��Knf�ն�XF��d�`V�?]�*(6Uhv��]���}�|i�\	�i�T� W��μ�7iV�7ϨS�^�#Pa�u� �hw���k�� ��[5��Pb�ih���\�;�(b����ם��6�Vk0X���v��=ϲ��=��ٜ5�����[D�D�!������j�K�o��UK�C"�!b�%�t66&y�Ou�xe�yG�Q��*h$�(�	p&Ě�;x6o$	��TO�6�߆9��c�:n�k������vƨ���ziS�IL�w9�v'����&�z9�9��s^�%�aQ�5W�TC���tn�]�E�b=��O���fX0����U���W^�|�ΰ�������c���oy���������!��Y#%E}xl�<���>�iP����q�$�U��H������.��E�C��p���N��%Z���r��ӯZ]��T�J���T�U����H��T����dc�t��?��ls=�
՚��f?\̼p�+#7�Ů�j��x�1����ñ���)t��M֤��m�F�������� � ��L�.��20a&�NU�X�c�J�Qy�|��L&h�#A1_���&92[�el���դ�r�I�^����n�e]��M%�:vw.�f��^����a���f�$9j=��Ma��B�9�e��D>�*�\��֖c�^�SFBQIA��#u3R,�Q8��ݻ�Kl{c��s�����}Ēiu�?���[m��<�n�[/4������}�+���0�u�ԑX5l���M��w ���0���B��U�c���jGY����,>9�H�=iq�Z���+%�ý�䓡��u@�G����[�k��f�I�uO֊�.�Dk'[�L�λ4�� Kָ2�L��ِ1>�c��&��-��2���P�=E8	n��p(�3-6�Ê�6p�����H���e�l���*��O�������e��K���c�%�e�b��5Z�{D(�R"��y|���(�/��ƒOf���Ŝ|ѧ84�*�]T�&�՚��5�w�n�����,���Cԅ�\�-`&g���3��`'���_י�ڋha��&x�5a��~W��v�F�o��m�qS@��l�m'�>Q�<!��-Ku�Ye���"��<�{Q��Jν}`fQHL�+��Ot����o����^���$�p4�!t�D�	m���3l/��^��!������F/y���E}�WC�0K����Q+�ob��7���ܠ�2k�
z褼�e;1r�<�o�g���$�C����P�n�u������MUsI����?̨�i�~ݙ[�p-R���H%�D�p�{m񆁰~�3�!y�0�����a�]M����`�#�]we�\�"O�G�r��'E2j"/@�IF���Ǘ���uʄ�^% 2��/�����y�!�<<��O�T[���U���f�$�9��p��ʯ�j���M�Ƒ��zQz��`��p��r�!�J��lVegI$>V��{$ �R��V+ �k�"�"�_� O���!b7y��끳E�||y��"�g�a�D�O��2�mh
(�΁���pQ;�[����/�����Ypb�,'��$���=,p�y��`:������JK��8hP�8;���e���V#�	�C���K+~K�����_í���,�f�2�=���hT�r�bdb1B�æ���ԳP�j��Ř#��C������X�Y~�`�H�\?˫�H�t��Z3��h����hD��6[-yk�5f�5Fq\tN>�(׷���XLH�&�>�;�4�5�k�y�Ј��!�T����c@��X�=�wXe�>�Y$�=�����oߟ>]�n�⡙��|,'����H?r�6��2xm/��4���u�KT$NAF��<���&��ۉ�H��9�К�u�g�'X��R5kc��Oz�O����1KL9"P��{��F��K��/;�"����p��k��K�
q�L�;ȉ]rFFo�i˚�od����(U���rPw4/!s�Q��)���I�	3�H��$X&�I�(M�������CA~aJ� �̮O���.7���j�`A�x�/�z�ЎAm���i�X�/R�Lg�4�g���E��Y�3_&�?`��&$`{�#I�=>���*f�Sh-�aG-8=0DrN?�7�pQ#�r�<q��p�[��:Ϥ�G+6������k?���|bB��Uդ���GD`<�1ǝˬ�3V=���	DF~����(ԋL%Л\�w] rN{c���k�0�FX�����_�r�����D��+�5��"iv�N�2W�'�����{�#�7�B��z�zţ�>۱cJR�/;בky�\�$ ��{����5���rR�Q���75%��Ol�'����9"?�8.�[7���OyͰmհ��Җ�C5�8:jsY��>[�@��Fy��^W���':����C���_��7�����ʢ`Xq�~tQ"O��7V�N��C��8�Q+�����E��\ElW�o�e�<%�=�;$��5+��S�=��hQ:V]b=+@W����Ok2̀��`�Xԋ���K[}�ڛTUk��[�\�}9�M7]�Yx �D?+XK�~��?8����*(�F�� �CQ
�&��+"�8��.��t�<������Wy(�V��&~)�4�T?%��\d��^+����R5�P$�����9Ѡh>i��X�����Q#V�������U�M����MQ~�U�[����֏����9�����-�V��!ϵ1�:H=�k��^9����2�BX<Yő�uz{�F�]�ő�`޾2@.��HUD�-�΁'��N�j�H6�9{GWҾ���/++9�4�}�FM�^�����n`d���
}��C��y�S&U>�n�z�{^�8w�������>�'��Vc���"� ͔ئ&�:��L���iɜ�Ho����I�� HN��i�/�?p��ֳ�o�B��D�)����>-�{�Z��ĘZ8�<�T�%A�S��r�H�Ă�rn9@���v>1R�+��C��r��ԍn�	�W�s���i�ݪ=����cY���e����HS��4I����H�����Pӆ9������^�{b��{�,X1tg]��-Iʦ{QWX��mo����$�*d���O}�L,gj(�Im���MU�ώP@#��dU�~a�^F�I5�>.�����g�-�JQ�~�7��}�4S���6z��������}As~兟�h%m���rJ�1ع�"R�)�BC�l�7	�M��U�Z��=\j� ��lu���;�L7x�0g�4�#
�mq~{Ws1��>�qz6�!e"Ekl��a�ġZz���qŀ r���j�W���QK�/!>xn�a��[I���楛]ѬW2�-�g�y�g�2�m�������Af�D$l�/xd���{|ÿT���a�Wz�ga�%{�@��Q�y��Ͳti�&ݡ �'k�4�}��@���(o�j3/�hյq̧��p�A
��+lsc�P����F
,����jM�~�({�Nم��F��S�]cט��RN�	x��?�Vz�o�\��M�nL�V����Nn.��A`��?�RƘ�ܱ�q�e)4vs�G4�j�����4{G�N]zD�Ї��)���k�40���,��V���Y�Gk�	|x�؉�L\��������b��&3��9&5�gh�rǵo'+f�r �zfUI\\e�8|��3���>�+2���֩���]��YB=b�c��gld�8��$N+	؂�=�knp�ޫ:\:&���-��e7�r��xω�"1����R1Ȼ���q"8�� ��hlT��#;8!]4~fJ4���3yѳDv�����F� 2v<���j�]�p�B��4k�����������ֿ�t��r������;�0<^u�
�����a��L�{r>�����܀�MDſ�F=(b*-:O�9 � T\�w`1�)=���N�B'�M�+`<�7�[��k���c�צ�z%zM��Ƭ}�W�@�) �}a���ь�ȏ��W9ƙ����X������A4l��Ԥ�W� ���'�1�- ^gP����by�>T�<����zo��w#�9|P]��τ�,;]���c_^��[�)RKګ]�J+�$��ԇ�!nӝ����� ���� ����R(�hD�SK��2�)��>Y�.�b��ѹ_e#��6����x��s�d�G��R��������̺hS�
��yF-�����w��Q�C�N+K�j�a�7k�1$���̫|�;�Z��o�� HG���je5SA�SI�؆��������(�"t?��$[��?�C�W\��U� �������^L�h���Kt�O,
�m{��w�,�
�0k�Y;�Z�w���Y|�$��T�̣�9���D�*L�2��Y�3�|������q
���N4��Z����'R�c��Nӂ���j����q|��F�M�3���8��"1I=SnzU����vi�(��'�Xި�R@�3��k/�X���hx��;��N�eQ��p�	�^k�x֥㫷ˊ5ɀ�&��t*Ɲ��ˤ�P������+�A������e�:2М�^�v$�^��k^��o�b�q=�����<*(�f��6QQ��[��?1�������ӣt��OG�=���������s��+'x�D�t�@�Ƙ@���WJ�z-Mo��Wy��(G�+�~�lA"�� ���sʞh�;5f���.@�qr#�zl�n�H��h�����=�,X�S,�b������E4�X���Qrb���K�/u7�p�7q� <A����X(Q����SVu�%C���F�x��:�7P����-��u=�g*M)�&�zN��4�H��$"�Q�l��C��6$J�1�j-�1$aW�{�D(�^W�ك�����4�ˍB�{���w:�O�������t.	5L�Ώ�yL:�EF.��Ϩ1f��=��W���_� 	%�=�÷c���o&��w�c��:�DE�mj�b�8*j�ɽ��L�&ɢ��0X��qH����j�cN��>%����x���M۪��� �W�4$����,�����{ +/��La幍�r����$�D������_���*�����%Y���}�H��8�D��^	T��g�}>jQ�7#�%��Z�a�/������;e�#h�Hjgg^��N���qX���r��02��hu�
1�.$��UdI�Ѭ��d=YL��8$�{����N��< �2�ok?�O��ԍ�)�X� �-vX>Ԕ����	�IK���"{����JK@�j�.UZi�\��WW����Y�5�޽�����ø�#�WoJ/�߼(��F�����PǙ�Fd��!u���3�410������N�����&3񔔜K�Uh��t�[N_E�+����`�Q��N��p"���n�~����#GY0������'� $5�VX���D���fG�Aͮ�C�J�t#x�7i�٠P���������f-���G���)d��Ӷ��`�b��8�9��|m1� �(���G��蝮��ov�q��D!�aC0h.ó��P(�K����]tIRjT6��l}�f5��j�M~IE5��"t�����C�d'M,��Cn�i<���wu~�u��bQ����z�Λ�LSϵ�kP�zrN�&bǆh��y���ʓЀ�����T#�Ajc$Cײ3�V3O�B�����!L��{s�_�7���*���m]�i�s�+����
"�������F���#����7)dqꪓ�rGp�<����nla<���	U}�<\'b��"�!��N̆�
$WC��+d���@;�	�ov_�R���#	4d�(��,�ٿ��k/��E��^CR�M���ZCO���9��-�;$��_�L�0����eH����#D/x����!F����W�<5K[3�i�d�=\�L}��8���'J-�g<�ƄR�ULnF��j�(�ZS}Ŀ*�'��~�H��5���~��p �/Ν�d�P+k0O����M��a���|�Iu�s�����}�cѢ,�T<k�~��zS��Nu��h��-�)��-!���$�}���9��6��g���J1����4k�-;l��;֕A����#	�*�w6���A����f����f}X��.��?e�\�'�O� ��a������w�����A��(5k���u�@9S�T^y��|Ȓ���=j�"d�L���j`'s��(7/�m�Ԫ��u�>I���#��������ߺ�7m�ɐ����d�s��'��b�O]��^��;��C�vj$C	&|.�	�=Y\X�Ē8��� g�G�(r�Jo�aVҴ�)�-��B�?�V��������&5.�k�������V!HW��6Kte��,�(~�E!o+|��
�$�����1�y�tg�x��iڵɻ��8�b,��=U�>�g�;��C�:���٦Jo(�똨"�%�3�M����Wrߴ��pb�"#4��4�����C�t5&��"B#��}������n��*(�J>��[�;��͙T@g��R�hBᘶ�쏈(�iS�M ��[Z�-k
-EIb~�?a��`��qXLpl��]�jS���X2r�~�2����,�T�;�lV�9�i��g�嵴��:�����K�� <�w|Wf�5��T�2��r1�|�~<q���o��]��)P��䖄��SgBS�)�Vف���AsT��[��/����<����(DU-))�:*�Aޞ5aH$l�5�d�Z����I��dCA�&#Rި+����x�wo��� ��3�y����{@����^�@����"%���Ee/,�z�B����l�ʹW��9?��8�Y7�T�(��v+l���<Wf£�|���w�/��fô�/����N�,w{�
��Ř�`�ΣA_�\�$��0��d�x�ւ2N�;щi�qpbB>=���L�2���N�d{�<yX-(C����&���7�Zw>����fK
_L��^2�*l�U��C�����\X��E�r�6�$�P�?��{�v�ۓ�pэ��3�	���?x�j���e�ml�2�Jh�vɈi	�}a_d�z�f՟bG�%c�%�V�2x�3�BI�1~P��� ����~�׵(��t��N=����J>��L;�vU�)1�I��K�o�Ȏ��P�Q{�y��D�6��/��]|�3ۋ���Z��@pV�/K6�
���x�
`�����.�?_A��Q�	�/�4���{~��b��Ndy�I��A��8���MI@_$+�xP�����]G�y�zݵ�;y�L��ʚDC��Pz�T)���x�|�{�)cA�G!G�:��+��٤d=��5"���E�'�ߛ��|+:;4&]��@���Q0�t�չ:��Jm��퇸���ү�V��~=h7�zd.ɹ0-������`ֻ�OqrƩ����]����T?�����R���A���˕�u&
ףN�ؚ��r�����^�N F��km#� �)HC3��~��bP%��o턷��~+�N���
5D��i��"��s�t}�{Q&�ܒߜ0b�ek� g��O�0P�������]��I�m/�,�{iNW�˼E-�0�:F����n��x�H�Z-���ɳhq��!v�>�Ʉ x������怏�w����K�Z���}�pey�f̢���Vl�@���)�ٯ^�˼!ݻ�<�xYb��4ѓ�D=b2	�VW���)NFZNy��ϱ���Tpq�C8�P1��R>��n�lP����'nNa���B�luN;ڧ���`��LQ�)����_@�n?�4l�%Z�Y1��;)z���+H�|�w�Z�����6�n�U~��q"�N�,w�2E��xA�G�вn���s���FF�	J��_�z�[n_�����h��� �����S�jz�UH�5k���a��7�x5F�K<��<����e��8�c�1�XChs���I�0>ZE�Gi��]��~Rt�ຣ���DK�`��� ���:v�"cDË@����v��Y��%G|��>�8{o���IKK��|��w���q^̇�<4�����Z�^��E��5SEetVIs��x
,�+��%$)^&}
�Ϝ�5�,O����<���p�bNjO@�M�J�v��Q����c��j�؃��ݚ�������؂���Z&�\�=S|��� �bh��t���(��h8>��~h��%�u?N{�Ny�?%,�ZH�d����=}�����SgY��#2�ԯM.{NPM���!���Dj�o��1�/		�mA���5��.�1<g(���9��ת#���׿CH��Ehz=d�Ć��c�Ml�%�t��8E�2O+ jsC��W�s�-f�+V���AWr��̡�K�a�����\¡l�z��p�u/����:η�	����Ϲ%|��L>��J�'��y��PG��<�j�N$3Ǎ�t$�6ߛ]<�������k�`�ZSU�K��u(Y���ъ�^��_���$�%�,�	̇Dׯ����ɖgz��������8Hܑ�]������BE�i�46V���XW�|q"��k�Exԡ;N?����C�ᚅ��ȏ�:�%��Xy;h�(����+���� �ƪ��4V��+0V�Z� j]��Nm��Nu1>7�6��vx'��V���\��-�3�Z�ۘ�	��4%"����z�SO< R0�W�3������@�i�Ϸ�l%�����2�}����F&�����c��s�>�Y�O�H�6AdB>�B�?��ݚ�T���>�Ko���E����ЂbW�\ۊ'p	���^v��� ���ӧU�?����ȏ�X�=u O��I�#c�:���UϳW�0��Ɠ��rp3�U��G!35K���_���*,}�j1�t,6=67N���<���"�!v��C���(�zځ:�;m(],jՖ�PS�Cd{����C�K̢���0R�&i1.F5L� K �q�rt�	$2~=;𴿠��'�PC�|S�wc~���G%����X�����q��w�d���!��+`���bQٱ!��R�i_�{1mB4��;=^�X`�+O��v��.D�@4��b�/Wh�q	���A����Ř'9�H�K�Т�H^�~���a�l�mm�����X�/93���$|�dcJ�і˅*��í�u��f���2�)��V%w��Q%�az$[��ֶD�Ȫ�e".8��-|�k�Cs�iU���br�î2�[Vw�{�㆘T$q��Gm@�)�Y(�2����,H��Y����m��i$\h"D
Ō^��Ǎ#��s<g1����|ypk��l@A%緳m�Y^꫋��|A���P�3�lg�n�u�v���Ά2ޮ-����~U��״�l�����A�y\���[!M���;Q�ѡ�3uoý�9-^j:�}+���R��=�P��,?�打�g$��]����A������@�."�S���bxzǕ���#�)Q:�CGa�?5%QU��aS'��j!���$�I��vV���0���D8��l�#�ŧ���˷ӈ��� ���|B��ʐ2�6�T�;�٢e�[Ҿq�8Kǹ���#̤��^�?6�o��E��j�\��u�M;�C![B>	g��ԕ'=��ʫ�3�pئ�؜�]�����t����r5>�CM�ͪS�� e��۟i	���t*�?l��2�Y�}��z�Bpʃ���(��@����p)4�ˢ��?�C�Y�Wd~�L�7ʰ�!}/�I�2v�_�2.F-�i��O�pl#,r|5��;��ʩQIzY��8ϋX���[��
�Z	���ZV����-Ԗg9ғqe/GV�p��ԃ9�x^@��n�᛾����B����=��b��4�#���&��l�*>��'���.\�/;��	A��He�����&������N�K���Olkx�`]Fw�-E;��_���}��~ S%�m5ȜY�q	f��Ⳙ3;>k�/�2:WD�GY��\_�R�(����B=�0�	�
Y��`�fX���L_@�=N�P�޸9�!�D[̢�Tp������(��Эe𪞢(��[���VҞ��x��(�N�010�<aeL���:����fT�|�fV��;�1�!�j�ح^|��R�Z�˶#�\����X��-4ŧ��c�\|�t���+�M��1�6{��uF)�h\A�����b&�Q�cB�fbz,�Oxz�n�u����m�]�80ӥKo:~����e_�|����_�g��������oV�����#K9�Sn��Ϩ��wB��+�4\�T	�_�?�mRr0j^�
�c�|��^�{��hMb���G������Jԟ��x�D����$��@�2Z���F�z�&
��w:b��5"���Q�h�V��g��u�ɝ���y%LC?�0֮�e�7��g�ըxzꙈ�/� 
UyΈ�n۲�ƍ�l�q�eԹ#�A��8��g����9�l�A	�U�=�8�}��׍Qc����4?0��"��׋�>k���c[�����F�
���Q�PU�(�w�aK$�ťu)�8s�m뗧�[6���������i9�B7����u�z�lwM��_�Qf�H������Ёit0Ř�97N2�O�f��-�.�i�o�Z�|��b�S��;!��;mb�Y͒)2�DT�����Z��Ny�E��u��wC`4�O$��r�kU����5�I*��8�	�!ػ2���k�i�O��*1�Ū���JE�f�._����"K(ǝDl~:?d�N��C�aC�|e��;�7���	\�u�1���pL�W���(%�� �c$���u�&DKhōjM��r5�>��I�n���$��V�B����L�}�Z������s���l���������Ԥ�+JNu��o��\������AB����kcÔ�@��8��!�����{�B�i�oq��ou�B�mF�(ɷ��̠�p�B3����OR#�4� O�S����R.j����}�g"�2��[4d筓�Ku��� �S����p��|��ͭ��^�PE���$`�%blf���$�>�*z��3�2��w��
|c�R�9�i��teD;Wer��컴�:�*Ak!�^�����Zy!@d�?���+�����������@3�-�0��UF�R�������ଐ��!�r?Q�ucyU�-<z�Sjv�����b�	�Rz�x#��_��� �k��������\�꺁��U9CFhS# �����􏡲�@����_�Y{���Gmg>��U�Yi�N�PG$����e ���aQBn*�L/_�v4���.�CTg�h��ƭ�����f�[�P���pm����WK7`y
y��ԫf2Lep��V��$�,���&%Z�� �0�?ob���|�%>�|�F����`q>>/���ag��߷���"��
 �W����L�9C4R�s�t�m��RM����fL��+vS����'�}l�(�ɭ!.�*����c��m�r6�������p�p���в�\�����A������-��Қ�i��"�2�p}WN�c�g�����F�6�B~Sua�;�Lͦ��3���?g��(�z3I�6wh0jk�F�a��4�n��v�bD�~��R�R�$�t4�"�Yti�Bu8��n����M�_6�uB�h�~���Jt�� 6���bI������K�t��?��W�W�ק�ʫF��ʳ7l���
����GS��Vr���t�&�\�o�.͛m�x�`�mw��VG��/�ܗ��ٖ�q�0�~;�����5���*2�~&�O����Q�.�Oq�F�g;�����N�(�!�LK�;����K(0��R7S�I��|m"��[h���m�N�{Cյ.@�j���D������lŗyd�]\R_��z7��/���c�[&��ď=�9����IY�$(�I���jR��u6�g%C����;X��0�4��i*-��y��4����{G���k���dM���Lw&0v�y3��x]ĩ4�����m��O*P�CV��c5t�j_@o5���u�oc�E�� �z���1gi@"r�	pG68ե��3 D��1zO^ѓ� ���j��j��C^��Xۅ�˄t�F:��)�0*��7
�	�+:
[fA�z�� �o��ey?�4nSWǚ�S?�Y�w���!�R\�bz����/�G��ݳ�x�c�;����}QY��MNOjE����W����Z#	�.���Tx7F����#��*��,��.����bfH*l���k0�s���ޛe�^C_���^˼�e_Zq
��̺��vz���: �i
W���D�WP���R�n�?`��z�% ��J#GJ�9y���G��1�n(%e	�	}�SZ�Z�y���`�R!���Evr[=�``J��t���L]�a���?fwc���t��"@�-���$�U3uR�{y&|�F�f7%�_޼���/��w�$�'w�]�4�6����<w*2�9���!���\�Ua���H}$�`=�T���F9`i�00�$987'�fbq�
q7(�t��~@u%D��6��OL|�e>PVG�GRc���k��J�w�b9e��q��>1�n�>�Y�8�T���\7�N�*�����<^����X��[�s?�:,��lf��ہ+��[���#I�	�773}L̛���V�	����Y�g�&&_�8P'l����w����y���y�@���LW�\X�u��E� RA��D�H$�f9NC���H��ɡfY��e��j;�Z7��ꌕ:����s�:����C	�陘���[Cp�A����=qЌKom��Z)���Y�+t䝯tH���i֐%��2�b���1�R�AÆ��a�|�
H��4���W(��o�����R&(�5�`�m���K��ذ�{t��@��ug��'����+k��Z�l� o�Z�ܧMPRKC ,)r�,�}�\�E�ቡ�p��Ѩ���*�J��Y1mW �!��������.��<͒u��P�#pǸ���N��T�t{��e�2�[T�⤍��۶�(�A8d�ۉ�S@lr��_UM��2]�<��19쎵׉�{�_k%��g/��{&���`\�{-~��?H$�����GR�`��.�Q�t�I�s����#68�S���~՝	#�E�|��[�:^-�Tij 3k���;w�C��:�7��G�)�2�Q :w�uu~�ޛ�8�,W����>�F$��d�ׁ�k�9�O�6 7���|zD�/�*g�Z�g�+���6B���EQy��
��2��' ���S�U<�:��L����B��	U	���G]��Aޯv�6�����893�aLy��K}BcTڣĄ��$wq��{���g�̀�vI�P�lA��^F�$�� 8���$4�G���M�f)4�-�J3'w_!��9�Pۥ�$Z1�@X�Ԟ���ל��" ����p;���10ک����"��\,M9tF�Ѫ�����[|q��D���	!S����#c���-�ٔ�!0�Is[(.��|ی����j�H�@N�����,��r����B:�)jVu}���9(�i^�U�>)�8����� M�=����ʆ�#:4�����J�|��fiĹy.�8�+D�g���I�z�1�Ό��TJ�E�J$�E��|ش�7���-Ȯ�\;֭�}{sL���m�>�M^��n%\B�I&�KA9t��B����O5j��@�h���W��K��������Z��=�YvUO�l6�^�c�J6�����mp��=�C������vkl;��NA'�q6�w���D��e�b��[���ZA�xVmI�����|aEL���ѽ�H�'��N�_��$K���8�1r}0XB�g��R`���d���/�%$�Y^5/�1 M�=�ܰ�

]w◾��R�~K���+��1�8�ҝ�Ҳn�7-��q�6��C�QgR\ ��!�?�r�%G`��	��\�
���-�b��Nw2Ԥ�ɉ���c�U+wB``��Y���L�V&�y^*Ɵ&z�:JP6T�K�D��ALWw9SN(��$g9�g�h7�yA7-�f�G�$��D7��ô5ƽE����-R:�7�ga9{l( ��/ʆ�t��4j�5�S��Kf$�NXJ��k��샐'T�Izk�Ò�ag��j���_��q'�44*Z�uȜ�E�:LO2��tv�5T*����]��ld���x�(_M� b�km% ~�L��z2�
�Ys�A��X��R����01a����{w
u�"TD��sP��\�6����^=��R�m�.���SkX���!���-X���EZ�~q��|s8_� |߆`k�Z�O��j�j����SK��O����#�焫��)��@�&'�l�w
Y/0`���"�����{R�J�i�B��G4p�@T��a�0���r�\�M�Ǹ���0>z���P3�c��y��	�U��o5�͜��F�}H�*"H���q�ܕn���o��z��i��L|X%�G�����l[��b1�{�>Y+E���u&`�m ��?݈��~"�~Y
!���q>�Gu�"2�=�;<t,r��i ����u��5� 	��`��-��t�a�� ��4��%�?Ĵ�G���׷���)�C�}d?��O�VU�I��!��E�R]o8��Vp����<w��v���]a�b��Z=���G3B��7���� �P��6��π����u9�-��e#��F� Ƌ�ŉ�(Uۋ1�dw�J�3�)ae�NA���v\�+b�g�}��6����d�W;��^�<���.~X(�2�1n�.���~��2����n�^��k���s�<����z��O�a"cb�<QvE����0�4taC�!�H ��e��j.Qp��0�3���7�V:DD�T6��4�K�Y��q|'e�E�� �>�舫ˬؗ���`�	6����{��kb��K/��#��� �M�<Vi���yY�Ԣ��D��,�x���T�jLB6�DtFRƗĀ�k�:ѝ�O�۩�ݦ�Y�؀�2mq���s������W)�����5�E����3���Q����bW	ɥ��2���xmvS(LI4��|�v����{3=�宗�ߤ>��V�Ħ���6�q;o{�m6�M����I�Ъ���ħ�-��oO��+�5��Kީ2|w�������O�%s�FG=Hרo`�!�uʿ,G�Szt��%ˣ����B���&�95�v�^��UD|���r�K?�L�c��JN11\:�-��Æ�8T����1 ��Vr�h��.�#I�2XP���E�U�������מ��_��+��	F>�s�қ~O��F�.^;��dB�:��ĩ���Ѫ�{p��V��`ބ�g�%���=x�O�Ys��]%#��aG�7�'�~is'oq�,�E�|���5=�^"�e�k]��v:&�ԀƆ){�93*I���)6�y�a�#�C�>2pWyEѺU�a崰�M��#����*9���Jy{�NG�EH�,ln�^	 Ȉ`�r���M���w����o[ ��L���O-�G�NG^T��8q��N
ct�W�/P����myL��}ឌ^�갶o��n���!�c�;�"��s�7ݒ��E.�"!Qӓ���'�!�AHS�y8c�0�Rx����q��fpsCڃ�x.-��4����!FeS�٨D�C���K&�b@�?�?�im!���<Zo ���3l�g��fּ$w�����ّ���3�<֧����;��`���
����w�0��\��(pO��ԩ֏?l�������c?��N���[bIمkRB|�za�Y�5��K�
.�,����m���<�i��è���#Y(X��N�
��̯�D"�EO:�څn�	y7��-���=����]==�~�ґ�KLǯ��@6�fqlwB��&t�D=j��Jg���%Y��͒���_�~	�U��9U �08�h*�Q5��J�������wٸMm�Js#������3Gv���\����ʑ�=�N4J�����y��;�ċ�9��Nc3��×����Og�F�n�Ȣ�ի����<�`�\�����n�������N&����i-�����3�xz�j�D`�z(h��LK�����28L��9�3ū~�c8.�>����ұ�L�W~`���h�zS��"�3����v;w9�����qwr�<���X(��� ���Ϙ�����x&�:h�
�Y��/�a��U�Ckp�τ��]�yPFh�X1"a�e�l���)�u|.X.��J�ʏ{�*d��"K�_�QK��Q'A@q�ȓ)�*���
�s{����gA���ͤ�ܮ��V'K��E��Q'��������84��,et��C��Z�A�44��/��}��#Đ�f�i��j ���I Y�<�X����r�n�`Z���ζ7��9br�<��|�v�I
����oo?nӎ#�C���̒��Q����O@1�V3WS��,I�qM'��j��SB�		t����߿f��oHZx
���*��·[�������Ɨ�u,��?��'�F�T��<VڂI5��N�Y����2����\\�ZPC�اJ3@��ӄ5}p��$)O������m�v���3�h�̵��
��e�C%�Z3�|�x�Z�d*��C�c�ǃ�3�z�N��͗�7��]��*<��Ju�q$n#�m��N�!6�t�C6��ED�]�J�%ΙbzULf�!r�LR��2��L�?tX�P~C��v�lu�15�Q�j}D����yULK�h�zP��廚J�iW���Mg�&{�`S�y�^>���ПeO}m:ЭUHG �Ǜ]�� ����C;HqO���6���`��� �	O���O��q��+���uF���9 j�W��`�&���bA�멣yA׼�x��M儂��䴼:y�lc�d�N���C��=�����`'�-�>����@�s�7�V�ϦNu��	��v߸��/��}���j���`��NI�} e�h�a�Nܴ��+9�༜�ֽ�9I���~�f&�1-Y(*u��M0��ۿ̐�0������9�d�PC�s��_ƴ�Ok5�)�����&c�H�$�8(	���3LN�],[63��L�	�by��fA�p�X�I���p8��2��f$%n& �r��c�t�?sGNq�r� ����:� ��|�2��f!��N�4+ނRVm��1�������k��O˩���g�n������2s/M;��zSLj����9.��#um�{�h�Д����hK����|Naa*�9�Z^/U��1�s�5[�3�\�i|1y��!�Ya�����`\���Ry&���ܖ.r�@�f[�2������ៀ��0^D�l��tͭ�o8G]��7tC)|���E%a��X?�t Ə"j�h��L�I�xw�\���G�"�"���a6'[�	�>�y!���lFO�4:��Ȣ�0#W���<t���=Yex�Ѿ���͔_�;�ud��6P!@IF-��O����@�H�rV�I7���ߍ��b�n��*����$ϐ�z9He5�@Аı�?�5ՠw��7	����G �z3h�Ώ�I䐐�{9�S����(�������B'1O���r[xhT᠈=>)
(��{��{B��O��Ч�^DtcQ�+;�k��P�U����8E�x���8�9�8^."���{����߸�9P��LD��Y2�������1�_�iw�9B�1ZSRF�]u=����O8$����f5�{����7to��FR�Dg�����ym��|����#��T.bT��Qt�N���N��AU+��)��z꿓cA���~����(^�	`tGW���O�EE�U��q�|��ԱA�AJ��A�wv��@L��	p�g�b$�n$3�B�#��>���x�n������[��_>Ȅ�B% ]v������д���LX�eE��Z_�1Y9虓��C�{6y�����c�d�օ�B��QG��T�櫛����'E��n�?�t�0x̍�ԭߚ��ʏ�M�u��x:�L꽱�!�8�M����|�E�Ŧz��u�5G�ۺ��ų��}���a��խsN�������('M������q�IC{�߁�����lq�?�f�; �C���o���r�?����-�S]�����q�˗Ӽ��%��_�B��H�2Ř.,�A;�q�=�֤c,B
ZѪHtP�^�]�A�h"����[�-?�6��#4[��и\������N�M�I@Y���_F�k���(�#���ߡ]b�2�\K
GT0�G��ȨG���f����iv�p/D7��r�P�k�9�PV��$���<���h��L@�����qX�01���0���1�q컱�S�&1\��gO͸Mh�=Жt��jS�B}s��x�bŴ���&.8�MSV�&D���Vt����w�r(��3��ě�i�ԩ����0@���3(��t�F�hZ�Y�����ِ��#~m}٦U���%(��
��ECD1jނw���Z=�ȱ9�(A�2�}V1�o� �Iܸ
X�R�Gpif��JxB�������j�"�/~�g�38{�"3�R��Wh�`?��	���-�	I���#�G�>��7 \�i�vJ�m�.�f�w)�B%�� ���}�8���{�,�4,)�4����qz�����3����Q5y�g�}	�B{�c������R��G��O���6Q���C�K�H�k�X|LA�A�N�*_��s�%�MM �"#�D�; ^� �������H�?R�����9���[�%������(�n��⑄��I]�u7�c'nZz��A#\B%���'�.j9;�'T�xO�@~�$�2���kuxpq���;�ӹ�i��u[����B3-�����E�oE��WHT%�:u��f \/!7W9�s�%�ɵU���L�C�ra���n	Op��}K/M�f�>�ު4��������p·3I<����M݈��̑Q����s,n��-�轮V�Z1� �vjz4� V+L�s�Eu�ȂEK��ٵ%�}ذZ�+�D�6�N]v:�s44�ܵqJo�ԟ1�߼7D�mQ�2a<.3���.����)�{$���rh�-XC��o�xBh�
tAŀT�;��5z���WK��E6���h�M~`-O�(�z�7	�ӒA�C�����������v.�_u���W�Ffc���S�\SH��z�r<C�d��<A�#l��0�+Gb�|�xu� T�#� �k��[�%Yh4��;�@�"�8?�N��}e�d���iR��/ �4m ��ު��9|r�r�����Z\<K6��6��U.W>Ŵ,a��#�)�/���݊���$u}��*�rh)c%b}���8<�y���-�zNt�E���� �h8~�]R�.��:���֐���:�Ðt�pAb��-��ǏV����a\��(X�6n�Nȝ��!�S��ݿd�!��p��m�@?!����T�z�>q�7Ͳ�SK�p�a��[^�(V������^�p���9��>ϞR�j�XhnDj��`o�N�07K|6�n��>�|[~R�n<����>@#p:]�:� )\cMs��h�҆E�d#���J�@�����&�V&�	oBߝ�D���|N�Y�g�7<�RfB�ȓ 6���[�� �qW�~`�C�{d7�61���4n)�S�
�,���{{�r[Jk�&��?�$�l@�u$��bhL"�~�,J'��+�wȺ�*^��,���"�����yA�o�L�d�w��[�O*���N0W'+9��`]Tom�j��;H5%Gg%�BYl�Q�t[�YK�"p���|:��&�`y����vL����
�����DMH;i�RQ?y��1:����X�zP�vS��o��������혺Ģ�Y�T��b����R����S��%b2�C���+�ǵ�
Uk�	l�m��GV�,~�{�Ux�����J��mGu�H������Ͻ�'�N|����CFp\�x��O1�x�^��o�q#���
pJ�Y��TNt�jImz��I���96]���Fε�S�:���Z��l�{��	8�b��E��a�3q�@0L�,�BW�j;��dvv�#�։e�!U�%���w�[���p�b�Ʌ�9&��=y��U�j�]mQn�T�D�E�lR��Ҵ4TH�����,4�ðִ� -�����5�g��$�N����V8N��̵�\�����fL�ȅ��d3��@�s�BVw)��KD�e��G�5
��C�����z�d/FS�"�t����<w�*����B�[ |Ɍ���*;!IF�MK9Il�M�lF����޼���Ў�$""� ��Ҥx`�����*���ϡ��7�Y�Nl����C�:��M��P��oi�o���K��-��?�f(z�,4r��+ː�������x�*�7H^��Uե�ؾ*[Au��k���ȕ����ucrb
r�#����6G���1���ݷ��h␌˭z?�;2	�7��H)m� �8'ac�Yjɲsv�Q��hv�k%1&���w�U�k	���=�~H�;�J����W�%Տ�576�CP���A�2k|hz]�`�D��x�g�]�xnҀ@���`eF<�� 1������`p%�?#��j�AK^�AR����o�ף�G�x������ �d��u?}v(�Ml��`���(h��o=�%Myt���dB�ɳ(��~�]sTY\L���:� ���H��Q�L�� ���Y�kjc����&�N��
��{�RX�!��Ć�Qjpk��`uv�H��Kp��j/t�{�P�_`F�츿�
!+�L��Kx��]�b�M�����ҊpQ�hfv��,�K�mۇ�ݥ���d_)�,�S*���4P~�.�{߄"-�6�8��8����bhd!��S۰���ùi͟[����:$B9�z�wW:-$���r�k�"�c�;ma}�L��4�љ�H�?"qQ·)�Uk�3������d��[*�^�0���#2P�ѫ��Zq��2��
�(;wFنk2I'Zn�P�30��|���~H�!O ��$��N�ߣ�� �!�@3�s=iLK�b���z�ڣ���W��	iG�g	ig�fħǡ���w�e�HE>���fT��㓼u�v�wi�$Wl���|�e��¨��e&����M���qo+�j���#LXc������`7���� ���b�4��4PC5�S�������9Z�����"'��6�+h�ZbO�|X�gy,�S�խ��U�竘�{ڹ���'a|���,B��'QV�*
��͊�<�-�FG
�����H�1�[~�:�VI�uY��t+r����v��Yn�;AAr��w�� �@�������)MT����Gqm|`�
()�������D/��e���b�����>��#y�����+�H>ܲ06v1�k��Rp�aEf7&�d\�dXt�N[_��r�yT�p�ԌL�A��h4�i�˚�jxw�1�xqr�s�c���7�b~��{?����?IW0��Ubͥ���I�/�4h�o���;z*�E���������׉>`���+j���K�M~�n�k\����B�Kr��|e�
��g�w��|�$,������KM8�i�Oj_�A������11Q����_��*���Xr7��O1��nI���%k���vA܏�� ��S��l+�S�x�ȹ.Wd��np���yi�xj������me��
���z�%$$c�8 �㞞*zs*И�������ɢ�-k�->g�VA0��۟�!7+ؘd(W-�!�"�>�".~k��'<|X���(�w'i�у��Iz����C��W���l��/h#�l̙[�Yo��^�����V����~�FSJ���\צ�a
�p�\ŁI6ſ�&��M����'�Q���М{I�V���J��<$f�)[)7�k�WG��x�j���f�sܣ�{��Z�V��� JX��xd�YvÌa(G|>��@����A }�{~�sJ�����<���'<t�v�7���f����0��QR?�����}�g�>�0^�^�׮Xԍ?���r��_W�`ͦ�b���p�
�`T�U=�-���nB�o*	E-��P��Y���NT�A��AGf�d�d�JB�j�{�.�Q,@��֍��m���l�ɣ�s��N���B�7��R���Z�Z���ù��S�C:��/u/����?���������fnH�~`A(��U��'nz�>����1Z��E�<�fx�0$���?R[V��)ND)_��&�ԁ��d���&�0�u��B}x�sڦಫ��#��3�~�]y�]��Zm�J�4�sOi^h�»����&��ŉ3/�%���	7�g�i���u�6.o��F-]ݳ�F��g0����,�h��o_��E�F�GQ��Ғ����6h{���R:�lF˽��~|"��RR����~�ʨk��bZ��4��C�� ӳ�����',�PuH@��i����o��c�Z/��vtp�z���_��/��$��G�b�u���158�nP�'��_��M�����3X��k���n֟�=1�g;�E�=�������>/��c�o�����"Hy�5����Bo�S��g8K���+A�6	���M���A2,��\Z��%]^�c/��su�jcku��#G��Z��o����Y{�Br�~�Y��L�����6���̲���+���Z L���<����Rt���M+��p�N�v�Mʌ^e%f�K+>�5�k첋hz%}�!�Ÿ-�rO
��?���\F3�1
@��W�n�TY6���B, O4�1.��.x0�؄����<����R97h��ލ>�O<�j#�-���E��Q'��
<~
����~b�1~D5�3���!�|,j��
<t�Y*j�-llܢfisI~�Zh��,C�=W�W�⫦+C6����ha#�z�Hy�J��?�A#�xd����t�(c~l�����Y�E�(�'�W���x�'��ߛ.����\v�mpڗT���N���C�c�m�ƕ�*%ܓ�u�Jl?�O:�G�D����ȪOb�C���+t�5QD�p7F��nr�'t���7Y��d�a��+#
eѯ��ޮ��X�MX�w�>��Ԙ�-�����U�+���5� �ȂD\�±S�_J�"���cd�3�I��+�C�OC���%��Z�9I��?��C*���~���Qk�B���O�������L5|�\��A9hYY��SMMZz�s6y^.a�5�H����l��;�
=?mT�<0��X+9�$X
I46:Ն[�Qߜ��>�PX�U�F�K���(ʁzM]V��*{_^WX���(2����}(��o]�1;�Ӕ�.�Q�[ډ����2�Z����R�;�1��ʠSM6��io����A5
��®[�쾛�{����d�!PB���k��c`vO23x\{�&�ѥK���H@�2�
Q�(j8t�D�Sɞ#V�
Q�8}��f�^��g�����ð���׶�M����'�"�����y�(3"z���D�YV�k�PE��𾄹U;$�,�	�HY�����m8�b!^��d�����?��� �m�I�O6�h�:ػY��d(���=TkؤB89K��8�#ɞԳ����ǻQ�9e!X�����S��Gi<��+��S|�����qRcg��]��{D�d��;�|��]P��փ쎦����kR�_�`�S�d|c4� mO��$~�׮35a�d�BIQ�M��$UP(x� ���n@�Ҁ�B\{��29�(�~X�춤�RDS�̬���OC�/G=�N��2�ʉ���z�f��E.�G��⎶�+4ǚ�Θ\jW+�!�{'I���2,F�x:�?�!Y\�ua�)��TB� L�"8�Q���*��Q��Z����wG��2�Ֆ����+l����a�m���R���PA��+}|��J�2��<ś���:>�hliF�n(���ɤ�Yf41��8��bASj�lf�R��G�7���P�z��;��M�j��b�� �	�7rs/��\��Gdk���ق�T��\N�ü��f!)����C�� v�g���Y�®���M�m��2:lF���x��%@�k���L���P��c���c��߉t�a��a_uY�q�=t�2t8�E��;��R������e�������|�r#��6���O�t�����MK-�=|ֆ�#Bk����o/���g�W�M+J�
�j����jP�n\j>����� >���N�D[?�������վ�����L̶���7ZD^lJ< ��}��-���Z�
AQ�J�U�G�el��W�{�8�߀-w 7�f_>� ���_�Ī��zh�<^�Oѡ?x í�f8��-�����v�7F�᧼"�Gɳ���xa�w�����PS��37|.�Kq-�Bm��/ƣ�L	�AfEBK�N�w����K�Rɧ��jU�WJ������\��}��_W�{��B��ha�e�z�<m���#�U�J�oZ�F���8��d��"�+M���m�o5�$deLFdi��K���v�2�F�İ1w��`P�0�S�Pei�-�'�.��~\���$(�A��ƛ��J�����H�,Ƽ��,�_[�����o[Κ7�.I(a<ҩg��� ��O�]A�F�B����Nm�??,)6į8?^۠)�Nn��e�D�XUf�N)��.�ML)ooȣ�0� w���=D0=�vt��y�N��6���b#�\�%+ P�T\���6���j)L�U�-Q���\J
��lO(���A���U�R�n��3m}�͡7�\��m�-��⎂�iߣY�B�	�s-�rc��]��};�dH��K��(���ځ�4F���Xal�s:>��P,`?�ov}���T���*�t�0�R�1��,)p��ϰ4�)��"���>������xm�mHFÓRj�cj�Y/�)�U2�$B�{l�>T�\��˶b�����*pe1����.tP���/^C��� ���,���J������S�,�m��7.�*s�q�����ҷԾ>��Xj.Ռ�% ��U�d@�͋]C���:�$g����h�D��lC&L�}�R4^'��@T�#��,*�/q� �r��_�,�����AXf#��d6[�=Or��2S=PLy[6$��L|^ԑ�XmÑb`�nϭ��@��U� ��~?��V�,H�u��
wCR&�I/��A�����(�>.\��/.�}�ע�~�<��TO��O�,�D_G���j�z��
�+썫ơ��>��x c�{�>��J-��G�����m��Zc�B�Q�.�L��<
Q�4xY�=�q�нJ��nn�Y�w`�$[�TάUH������FՀT��;���0�u(����ph6(F�$x�;dqW�m�٘0��3F��ٶ�0bh]*��� �^��)]%0�*|��3���l�4�=z$�Vl�b@���58��_�3l�����;唹ބ�O��{68��O�ZM ���ݻ'R��S��������N�m.+�C��[���X��mH�/a�rg��l��M�_r� spǮz(b3z)NS���Zѯ��)�Z�Q�Oj����#�1|oɛ��r�&+���m[R�O��F	9�S�LN�m��V����,�i�jR���Y'��`�r�7��Ւ�6�f�L��b�%�̎�D%6$�	�n	��Q=P?��:(���t�K�����(]#�S�"��˴�U�s��އ~U
�1m�i�e�8w.�&��`���2e���z�V �Bi[τ�ģ��an�CDƚ����c�z���ʹx�a�yYWA*��C��È���{�3ؔ�tW� ��	�EI�O�í3��	�e4�XE3A'>~I�D����;2��Ⲿ!��[˅���Ϋ��+/6�r�e�\ն0�H[U�8���Rk�]\���3��q]��<._�^�|Bo���R�E�<�$B�GE{��p��o��6c�ț0%}��>�VH��̶|9��__~��'���k����.�#��&�j 9�1�hI1����������K�AM�tՂ�a
���|0,q�>(���$Te����T�^7�ɺ��S�k2���@������������LC#��c���f\��(��87�渉�^{�N��e�黻�Y�c���J6�ؑ���3[>��/�����X��8ǿ'����c<�	oUJk�Q#�鿝�\���zjx㎪��l p/9�G�G��1�� �Cub��zp\�u�os�{�M?0x�I,eK��R��C$��� ����î�>�8��z'�Ϲm��A7�I�1�&��f�����3����]���6�����`����˻<-8�f��������:��sXu2g֢�`��)�cf*Zo�����7����J3����m��{N�q4�m���}*�	Awd��E��/o��V��&���H�� ���%��C0B@e��R����|]Q#��k���{mAC�n�-��JԻ�1���6�T]e,46$`3~gB{ϼ2�Ng�`\4|�+�x"`� ��k�H`1���S��,$�(C����W�d�r�"B�h�@���%E��O4�E�W��!�ߖ�;0�>R������.���bV��^����v e#�P^+�H;X�2�˨�|Gl�W��% ^d�͡ҩ��a�>�*��������6�?�H�(C����]��O�.Oq�i�t�1�}&�Us8 �0�������,���BH� �0].�a�:M�)��HBpT��V�*�o�LQr��v����8�6�Ù�[y���Ti6a���i�ӂ���%�&@'T /���t�ף�Q0�ɝ�i����%}35��Sƞ�Cp#���@W���*��L݉[=T����9��3)����H�썖���g­�Xvi)#����$*��4-�OO��dB��+�6��O�ܯOcԧr�?i�\@��w(NJ����Dm��t��OZKۿ�z�¯�'?X�am�9�u���W�,@4=�t����>	� v�D��=Ff�o�)�����@<���ʏ��ڏl�s)�.��};=���ZK��H�(D�=~�X��b�[0
��BP="s��N�`���s�0:�>�.�v��H������@,'v�R}��4���s���c���>�b�v�'�2Y�5YbF�<�����y����N4vK_7pu�i \�s��
n�������t�����`��J�[�v5����l69R��@��V���ֈeP5�w�c�1��@����h��()�§T��ve�glW/����Y��Cv@y�����\��!�Xҥ��V�14�$!ލ�Nv|��l�jT�Fx�����\���zkvo)�Z$R�vp�+���Y���D�IdGS�+P �9�����9E�2�ӔV�fY&�N���g��צ�ԫ`B�8?����������M�K{gPvG����������	C�]��aԥ��יV���D�0���l�R,o�QK���F����	W8 �M�C�^�?"w>��勞��ؐ�D^�`
�L,�_$F��>p5��f����&�N�.!J��<�z	�Ĝ�vWy둬λ8�jp��Gq@���]ƴ��P�k�M�81z3��]���â+���Z'�-BHϰ�^t�i�a:���]�����U%!h��[��Zƞ''��Ll�T>��v�;�Q~�pf"f���Axp��è�m��l'j-��b���pX�L�c,�3����u�-�C
.��J�q!B��)��I�* e�b��ߕ��]�5b�k�t��H}�H��%'�T螺�Z>��~�2آ����|���+�ֺu�����L���$'��	��Z��<64[H���[�}��˵�{�2�O�Д��?�4�p�Fæ�����`ꙟ-+�8���n�Auџ^���/�Q�SG֞褲���$������^�l��>=�'ɸ�Q'�>�F_���_T�k�՟+D�kF�c�Do4��8_�
��W"_Zrq/{�Db`㠒�v�uV�0O��*�
��辴˜L��,V����oKa×=�6�����}躕�
)�1��$*x�x5)qʇN�9����!�4�c
�up��=�b׶���<��W��G4Xx�{��$rh)��9�%0�k�́jf�f9C�$A�k��(��f�D��Eud�)����b�~��ќ:qAR y7x4A�%5髭��_�Ki��j����鰓E�(�	w�Ӵq���Q���P���1�/zN.#l�!��r�i�`L��h�d�r+CX��;\����<��4�~90�$]�8%��
��zΑ-�O�MX
�n�$f/֝�Z�v>z�}�C�JP�f��ybƙu��SgG��銼i�I{XbU���~��˻�
t���h� �n}�f�Ȃ��3������Xݎ���>Ԧ������4�!�,���`�oƙ0y~�B���Sb���"�D,�1�1g,U�Z�v}��D4���JXw�I!ű�s�]gD_�w�0������j��c~�M�����V�~Yw���S����B��I>Ɛ$�-eQ��k�,��U��u�	�k�ð^u�yT��d�((df����	�yq�E��{�t_�n-��"�#0/t��hm��)���L���(Lt�����{`��c#�ǰ������F��F	p[�*!s �A1��Y��r���x�i�Y���_��>���%� �k���������r���m$Ze�jB������TR`�>��}̵.���eƼ����m5	E/�?K����լ�X�&��iC�%W׃�\���b�� �׌�ۉA���X�����a��h����iɠ���"���;=����;kbx�<ev�@T�t\��k��ӳ��!O%��fN
I{!=�7�� ʑ�O��k�6 \���|�d�k�u����z�	�&C*T�͏l�$��Bpn�$J� S��-�B�W�+V��WS�$��.Ȏo7�w����Q8k��$b��Ry^-��2:�v�i*�V"qVk��P��َ���<r�=�	��ն��8��ݓ�[E
������r���3�E�t�igH$:q�0s�&%��Z<q�s+��;nf�C&��������)x>/[�ݛ!�2 |1/�-x�Vf0���]箱�ΞL4���k7N�߲4���� T-��Hi<�V������ o�ɖ%��o�11d�B-'uW�E�]����]��d'�_{��/F��F�V��{HLKlc��m�~�^��?tM���s\(Udg}#��'bMݭL���Nn������*��T���k5K��N-��� ��|�� �N���$9�߾$�Ue�X�SF�#S>U@�P�Nz���!��6��r�L�g1�WdU�8u��H*�yò�
�Mny��/zT���=�+a�d%��vh��).d��C"���+<VTD��?�U�sFO�K�AFM�G�<�,��I���@���o�_���ڝ�t�5�z���G��C:Gq���Eva��O��&Bqt���#�^�����˸'��]�񼄁�u*b�*�윒Οj�ͤ��&��>��� ���_�썢��9̷��Y̓[r���Nw�:�[�ee,,���μ�:�p�FT*�fQ|�D���!��v���vN��@��P��g�|d-��v���Ҟk������_.��4�z%n��K�G�-G�	���[v�8����[ hs�2>����Ϛ��=k$�[K»�>ź��+W&�ѴÑ���k6������2�1��GY����Z�7�\��9��yoU�0���j��b�z���3�4e�'b~5�/8J��{�	�i�>l�	�
�J�.�W��j����mכHz.�UG��ad���K��H�J�����:�]����c�NC�q���2�F]�}����z�`��h���9��o^a��Khr/h�rhy�`����SjBY�k�ƙI�,��d4_~��B)U?�@�����?�#k5�C��9��h㐠ON�ܖ��}u�����%�Ф�3��t��k�L��q�{���j@e__+@Կ\�,�w���_}f��Tn�H��5�.�EW����I5'���ac�������;*�ߗ*@/��NY{v��q��R����{��J�g~;&��F�vɞ�U
~RM~����*I�����l�y{��L�g�:)�{4�^�Q�T���R�n����Ou�f�A��`���Q޷��c�?�"{ƍ�J1����@YX/JF�Uk�,��$�OM�#��D�R��C�@��i/kp�q�Y�p�ހ|a�Y�(g�'�D9��Y�}���в�:z�?����	�[����X�����_iJeҏpH�kL��s8�W� @9�P^����������5eg�:���o!h�/����^L/2��O\�)���s����c��.��I/Ҹ��c$YCϖ��9��4��5��p�<S4��a�Ʌ	�$�ex2���mD?(��{6�9f��S~sſ5�=�Z�=dw��v.jT�S�K�e(��O��ꥮ�\�%����By'�lŰ�U�^7����0|�%"聲$��/�ȇ�S\����b�;��`d>-�&���شmL�*U��>����l��J�h�'42�����)!�-*�腽��������4x�;�\[8�0M�q1�@�NTi��g-6z9`zzp<b`_�v_ �)?v\��A��#���qa��`SA�\y>W�8���7�## +���0��LV�N�=*����k��5$�6>[�����t'�Gb;05�
��F!��+8/UaO]��W��w��iۖ_ �n�(�O�dmk�\�[ ���c24_�I�����Y���[���gߵ�Z����A�#�۹t��kـ��sq��T��ϴD_�ژ�J�_� s��6_�1�.s�:9@�
_�P� `�3F�z)�/���e�q�9��c��j����f7�T�"�A<MK��2���1��M"���T����l��o�3�}m�L�*O��g����o,7ܰ�"_�m���&�F\�SQ%��2ӿ���0����ւP�������� ��蘆��撾Z�[�Qm����.&�6/�!W�̹�ŒeL�K1wH	�#��&h7��MC=0�h�X�����2���;`��:�]sD.��M��^5H��*��B�ֈR~�e�sȧ7S�4¸�K~ٻW}�����m9��<�y5��S���Z�>f��\2��?��K��x���?
h`|i��Dm�������:pl&Z�����Ԙ�ew��|pݹ���Ώg?	�'�s/���:��ިߦZ�K�]����=i 7��A~�v�l:�����
'b����[�!r�=4��b��� �N�Ã�a�i����bg�C��2vJ& �!�|y>ɸ~�;O��1%F1��\��Ayy��W�'Uc#[S�UQ��c��%��B����_\�A���!��W��KPέ���L�%�TA-L+�@��髥f# � *Q楒U���\�Oک�����@Gn��|�sm�?�.�}P��!�@�6͞�9Ʀ�b1>H�w/�_�%((�o��dF�ғ���13�a�o�ԓZ��,��hP=>I����
��WI���7�K��?��J3�t�mxH�s�#j��{����Z���]��,�l�#��C�X�HJ~L,��cJĎ��<�@E%��4D`����	�|)���L�S�ë��Ő&��߾L�Y��Dv�\�����!�Ĩ��j$"4_
	.r�R�� <F{��[M��/RQ���H3�v|7��`}|;�
Go`,\n֙�e�q%~/s���vX��}������^�҆��ru��XI�Ä�8���gF�@JYU=dPyvn<�{�n�CN��n~(�����E�}���G�g��N���")_0����>(��~S�n����_�	�5�aB1�D�k�즁u��4Á��1��:΃,���+��{boG|n�n�͹D&m�1&����u�tˣ�t��2���T�Z�]!�C8�h��`���.)����5��k��L.}����	!�tBX�o�%�YR��o^7�(��	>�xM�b����w ;�}�/�|s�Ԛ\�w���ɽ��}�=o j+�~�w]?���Rv���҃�����pR!���F��V��h}|ahZ���7�M�20��"8��w�S짭�=l	��4����k�O��d�X�ت$�a4ed�lT?I�\�S�ͯ� T�4`yܻ�&r���A���L��:?�5�<��$�I��a��j��ٚ�ܯs��W
����J�]�u~�?/�NW�#�����l�u����ϭ��ܟ�3�*���6������y\�I蒍���D�%�:U�XrwE�Rm�܂��u�pA��dsYɊ�L-5��q���l�I��zN�=��P>mB��M%��f�����K���h��K�U�n��+~kk6V���[Il(px�x�<&!W��W�z���)P�a�:Y�9�; �p	��-
K��/w�N�ZAÁ=?���S��^1����aΨq�oU�B����\��W
i���y�w��ϳlkd�à�d�@F�G�}�L��s��)��G܇Y �f�)��~j ܉�z9�o(�2��1;�n��c���*�>��K�E�jG�<���Y�28��AF=���c|�̿�}��t�ѓ$��Ҕ=�ɤW��_�hX>�����r�)vF�635n (Q���"�Hʖß������k��h=:bf��I�
1�9�N!u��*̉D�5}�]9"Mw��Qq���*���>��fqM� b��9F�|��.��x���4�Ț��3����W|@� "�cF��I�\6�E���,W���\�^�$t=�9���	<J��yRޅ^u]ܺ�W�"��[��gi{�^܁�E� $�|2�:�ꨅqE&�뼀���F1���w�2�[H�:+#�H/��PTT��C�G�mq�6JT0U�6���?m��^���8���>��2�{"H�P�X����?�߭e�?��9��$e	�~a&���E��â���0�mQ�<�=4�tzh<J�`�����E�0��'I~g�Q�R=X*�pS'�=bm^t�39���@��渢sM��c6��s;
Z�j����f��p�Q��H��dw2��ų܎���X���v����~�J�x����ēH�S�����'V���o���25L �c6
Ջk d�=8�:e,��Fɺ:�����B��9�C�Rl��O=�f���o� Dp	���D�S���5{s��Fv!���▎R���Д�}A��+�؀�dʲ0`͢'B���A�0�r�0�VX�=P"Jk�]ǐ��v��*JΆ}��-9�Bb*�
��j<��.LN#�#��,C�"=�c4��R�uAr�>���Q��2:%�KaTS}kv��	5�?p�9��\��_UwY`�H���s�G�������1{�*��RQިTws]���*ڑ+RԼŚl�m�X7��Uz.���_`��uj�|�L�ؗ����A��]C(�(��4�'��7��Y�L��d�������W\�g���,��R�e�� V\eU�Ok#` �-�- �c~�����ظ�k�w%[�� �C��4�Oa`�s���
k�4"�,j�Dد�<6Z��Q��X���6�+#��1���,���6aADZrTXffٷ��jegfى�)W�fٴ������,;������L<)���"��-Rd(�Iյ��ӊ[�|D`�����ϻo7S�<���^J>�]3���wi<w[Z`ze������'ƿ�q��(��?�G�^���K٫�7����Ŏ���x>@�b杹h*�n�!�_���L9Ƭ�O�)��`�̶y��e9�ﬅ���#�]���,Z@����\c[���?t��!��/=��{r-tF�Q�͂�Z�U���MsRP����8��$��u�|f���59)`V�ft�D�m�V�K��[�!��,d���0nX�!]>��O*dq��J7��O�����鸷1P\��q?����nd�9�[��<@Y��Z涳�! ��m�����>!]�6�p��->��*��M����ە$�"���)�l�.�-`+A�2�^�l�y�+ഺ����ߴ z�-�������V���I� .��Z�8�
�4���4X��1�x�9A�TuJG��v��-���d�f�y�d��b�6h��L��>`����Ta�:jӯ-FqГ�L�\h{��l�W�(Y���ɕ�.��=u��Z�V��Z��+�G�Ra�H�����9����#A��� 3�8sl�Z�|^m�H�-s�)�eaL�V͋Ϧ���F��C�e	ѽ �x�tfC��%i�t�>�Nm����.m̹$$����p��#�N�y�Fo�]s��%ӕ��g��!�r��a�eB:�h\r�ٛ�֌���C��k���b�[�6�GS|YV&k�:����*�}�~K�ʖC��O�4���V�?��������-5[��Wom6�4wd#���m���u��5�����bQ�x�"�,�';��[m	���Z��	���Q��PI�qj��K�;Ƨ��׳�������H����hl���ME
����[k��Cɬ
Lu�0�L�N�SE�Ώs�3����vX&=� ��:̡kA������R�(蟧c�ϖ�H���\E�����7�����E�Cw�[� ���x�w� �X�E�����g��i�jSk�Ɲ��w��3?I�],���k�Gu�c��9^K���j?������-D`��L[���`j���Y�J�������֭��Ɵ�ך��bJ�ᆏ�v߈�1w7���uK{�'��[9���		>��v���n�B����`} ����P
�o-(Ne\��*xW�;�!�-�tn��@ʒ�	�-�J�����(p�.@���8�"�#�f3H�@EV+�:T����R�+r�Dkd�J�&�Y%�ྯ�������1�5�]��GM9�07�uVԁx��u�h�[q�կ�x�֐z�1)��:��C���Bȥ�8A�`�C�wp%���c��T����6���ϫ����(���;w�M򔃄������jW�����E�����v���	��K���}��~߾��zLL�&.��	 hQ���s�9��������2z��+įg�h�������J�)�O*�nDm�fsѬ�~�Y�\�a�����FK�U�i5ձ`ND����8���1���J�����#x��i���n��k�ޒ{��A��X�x�(u�oːr���� �5x�1�rw��d���>	u�܍v���k�ו�����R{�#it)}䝻,m�̝$h� 1w�'
�A9t���
����3=v�r,�ׁC&}�t�?~Ad\M�O �	�\\t���^[F�v���ʃ���\��\�����aФ�5�b��qP�����ݪ�eI�Ws�t�5�	ӿ4F���Ŋ
�W =^������6RԪ�%�(����߷V
��m�M[�&�/�����/���,p��u����Fdkr+�J�U��CKY"� 7�|�C�$q�Iv�D���.�6+���/�>A���\���Q��6���[S�����f'��]���]#w�>DчI3@j���@�pQ��q�iD��9����0�^A�����nn"��A"�n�����Q��1RЩ����b��CW��!i����1)QV+FN/΍�s��&%��2Qj�o�KX�7���ҵ���L�Xї����-n��y�ZP��0�Je�Q9xcj7|'���$����.\��n��_{srA��x�\��7'E�P�)�[�~�/A��֧�O��W6򗗍�ĉN����=u����:a�E��|n(xp�u��'f���5�O���5�W�-��O��R�$-��8�(YLh7Ӵ��O-'i��A�j�(���r�bI�5m�5�P�	f]�ç�M�)ރ
�O`��9s%o�����QY�//��,Ǯ�{z��Z�Z e�Hd&����
��a�m4���p ���S�|r,|�H_S��e]����B�8���L�o����~������Ix<�X2�B���AL�^ƶ飡c'�^<
$\N�1/c�e"`#�,z�:���{��==h�
Z�ӛ(��6�M�G�i�a� Ό��]�oQD������x����\#@������d�ݲ��B14��:mîԶ�
�����O�I�`����9��,�M�1I�*F����T��,4��GՏS����X�72lY�  ���G͘�m��̯P�]f���Hg�x����ٙ�B�B��` �H�>H)[�l_�|�����0$'�k��$T���{���)��Rԑ����/˭��(3��wC��X$h8;d�"!�_�aL�	�	o=�ў���*zކ���F�+r�nS�A��c��v>~G�4}���^z/�zMcX������o��л4bY4�EQ�!WC������"�����9�3�?>�¼��zI��aY���8Klt|1t�]؅�� H�i&����F�����|��8�\����ՙ��d`|�w���]�m2�XF�2l���#	�M ǉ��T���s\���7![>j��u턑�8���r
fy��jÎ���R�췻S����V��ԟDN����Ő��P�d�m�Qu7��R�<
\+��G9vR�'G�&�F�N��kJ�F��?h��	<?
BP�R�}W,�����u쑫��)~7C`�.tr/؏e�P�W�������j�Io���ix����:�w�{�����C�� 8���i1	S�cz P�c�T���i��'09�������a�O]�"J���^�q{�����S�Ǔe/T����ږ�3����N�&R^Q��t���W�nW�����Wc��Ũy,�s��L \�~�'��~��I	H�����J���щ����N�����8s7j�gs��%�2F�\�h5U��H��f /@���v>�VW���7e#���t�c!����?��j�|�gv����a�bX!��;��g̅-�َ�o%�hW��Yt�||�M�#�vqn�v+���M�Re�Ax7@�g�*�3 s���jǠ	�n���,+����K|1i%~w���%�>��=�Ԓ L��	�(������&�U�&S>�$)�mJ��SzTa[UhMÎ�]�{�O5*G>��^��H��50[ŁPX�$㽮�'��
��(od`=���_�l	L�U�����9`�pi���P�|���p�4B�8��:����[@�c�/|I���̋h���|�����K���ڲ�8^H�n�G���y�ޑ��Ǉ�ԡ�m���������#�BN�Y#�`-y?�� �Ȼn'�����	�ݸo���J�'�ek4e����Ku�>�ߪf���s6q ^�~&���ptU�:v��DP̾���C�Cˍ����|z�����ң�јL<晃&��e��v�|�>�w� � �\r^��
?�RUx�dj��u�9�f6�|����/v	���D�&�hq�g>��J0"�.v>"ҁq� ����T�Uk������m Ֆ��,
� ו7�G�V����Y���F�"}���&0�Ns�f@o�U���{����0L}Bw*@���q�E��_�z��8�J(�>S�P� |��ӯVĴ7~-_�b�C i ;F�J@(Ә!4R�3�(�5vx���YQ!L� y�)��w�2�d�]���$f6��p
�e��߯�h��rĠ�x�ɒ��ߎ$ƕ^`��w��uk����+�h6��R�w
�t$�E�0Rݿ�Lsûes�#^"]���V3s��o�d����i�3�]��a���dac���+�T��B!0y����)������g�Z��e��~��+�Q��t��[N�bj}�5�6	g�y^:>�&�u4�:���L��?T�x'��F�"���k��'Vb��O�V��qt��G��}yA���U�1k�PG�'.s]*Q1�t�lh�q��y@����Β]_j͠�/#��i� �ū��O[��<@: s&Q��>����	�cz��RT-D�F��p�-��PYeʦ��w�u�-�@~�;�7��:�1��x:��H��km��j8�p̲�������[��􈑃�j��#?`c���c��t���=ũ�o�@?��Bd��,{�1�H�_�}�v�_�b�G�P��3"�'E�;����iQ�ݒ���V��H�j�Q�����z��W=h!��l,����*>�ػ������ #��Į�T��F�9|D�]��Oｿ�{�`jV��Q���r|�byjMd5#//}���*y�gH��>���%��҅�%a��bl=��B��0�����T8#���`����!ԏ8[F�����f���M5g��I7d���E l��^�֯7�ƙ�H^L��_�ĕ 5��C9�6)�F�������֨�����{tj�m�&-��)`�8ZBh�1�kޮA �l�5���'`��e��/g)���R���<� &�s�a6��Z�X�Fx	[
�A;&�^`�ţ$O�����ӗD=8N�o�.�P%�6�@����*��M�)���:�!U3ús,�_�8�:����"O1�pT������"^16'���\�!����T��t�
�#�`�F.�^V�'|=��ߖl����RW4��C�Ξr6$�U�uq�Q��'m��o܅4Q�#7����������Fy��(/&A`m��ںO�E��~er�}�I�0V6�������+��zƟ	C���y�٤��x�:dĈ�i$}�3��]Oj�� 3��_�ٗ�������r�G;��g�V�5�K��g	���ef����=�� 'wJ�eʋ�����t��l���^�����HH��xO²'�
`�<�C@�c[K��2�2�/(�/�ۡ,�^M� hLâ�E_76UvE�!�M
,�]8��XT_���S'e�dY��u��4���e����wl����4$��0��oe\�QB�;�i���7@��z�_�]�� ='�k�2=����e�:r��L�*r]�*>|�`n��7�o�0n O�	w�A���&�9��hs�Vd�n���z��7�>䝲�F�-�y[�btB� "ƅU�X;���p��|Q�v���kZTF�t 
��_ �XϏs�d�"����Z��]�R���v����3�\<����}^V��%�D;���!���*��._�Jj�:�H V�T��"�7Z�<��ݥ�}�?<廬��'.qi2�c�
��)*p�L�I��0��,~���5�z�/����;t�% ����pz8f���Ϻߓ9�VA�ű��V���MqD`�������!�a���l�5ҥ� �H���ٌ�8�n��){���=��*x=�G:T�n��;�0�$���SU5��E���H��<bqW��y6��ܕ�V{��/F�� =[�U���0�;

� �6_Y�ߩ�����Fȼ{��~���O X��gt���.0��߇ۚw�o)�b�KKd��c�q�m��� �_�s+.��$M��\�Cx�V����{_&:��d��67��0��M�h�"d-2X��kɉ꾜�*�R­Zz�#���i��~]I��VϠs��b����*��#��?^�>��q����y�آFʃr�+]�My��˪d8��K��l�:ڨ��'���f��Nj(�m��,�[�){��M�R�$�\�5v}�FQ�H8E#����1�u�uF�ga�*�f�ܝ��5e؋+�D}�+{�P( �[#�v��cST �$��/�jQ�+�Ι�,�Qc�cyy#�J����i���R�%�(�<&���������(��3�ϔǿ�T-/�ϯ�ܾ��Ss��LyL�G8G�B��V�thUE�ȟ�`a}�\H@b"J�[����RT�`���~�7?/��#�.y��P*I\]]l~����VyԴ�Sx�&}}�������� �Fܔ�h�%�������7���+3s��?�5�΀J�$Ya�#��FF��&���A��e��aH�\ٞ���^�D�}H���Hny0k���u�Mz ��o�tJ��T/2�9U�t�?n�T��0�C���'�Ԍ�rm+��L�;�׵��������Fw�6?����qJ͘1z���l1�<F<|��N����x�U�l�.�cq�*��je
�\�Y�����]T&��7�lؖ�B�nښ�'�n�������(�Ck����益I�կ��C�Y�vY�$�j�J�G���WHy��1j ��[��k�f��!�1ѩM��73pG<�T���5�*�R�G{1�}�߼Lؤ��c�Zc,o_w�wɜv��cϰ��
݈à�e}��C0�ځ�P��	�s��{o�~��;�;I���C�Ok�������¥_7L�� �9h���7&u��M�pw72Ed��%�_���9v�ٶF=��a�D����u�8�&D	�pe@Y�k?� �\<{��M�,����]�2�gw\����{ ��vv�]�����$�pE�����
�0�N��f|2����_Z��M�a�J�3IU��w��qx!+1�&���^B�f�n�����T�����ٲ}���F�;�^
k����. D�}�Њ�t�v��i]��QSve��tݮ�hN�ݥ �-�Ɲgj�u	Jĵ��3V�&�q�H���8���i��Y�kYJǺ��Mܗ\3�o	�� ��wjb��a�=;o��{Y��񪫰Re����Ϊ��c[S⾛�MG��S\oW���D������衔�17w�aK�5��ݟ�Y�݃%ң�'����$<;pO���A���#i�	E��_��:[/[sx��ʺ�k�&��%�+��rd�a�:[(XsqGb]��O���9�Р}=z"N�g%�HY�E-�i�+ά�_lu�8����s3)�!�d�j�z�t]AF�J�b�GF[�T�F�茺@�ӅtלmN.m@E�f���L���=Zq�ޡQx��$iY+a����"+h�	/�,��h��_ۂ�Զ%��I����,Y�Չk��!����</}\D�����O�V����SQ2s&��نK���^��d�˫Eg�2F����g��y#����(��u�!%+���	�د�L�ț�k��
z̘�G����񦆼S���:�"/�&��#��F~��ˀ���C.���$�nOp��P��okW`���?� x
S׳�9���s�{2e�x�:]���};fDb`����&�q;J��N� �]�niš��A~���@m����z�0Zq��U%�����~�HwF�&!�V����M�g[[�J��P� ��^����k�0��N��/�@���"Ǉ�~�싔�r�P���%�d?�Nо`'߾��.)���͇�ݜ�!���o\��h�n鸞���H��.�� z��ڙZ;S�������"�w���|���/'��Ta�5��@Gp����4�sJ �)���νW#�/\���,.tC�����������ܖ���YP׃���p�"D��m���0ϡ�`��_`k��B0���4n��rf��=� �U���I��ei�
�n'` ��p���,>�^�Z'�a��#��a��y	G������/B��O>U?`�Eb���=~/�pAkgkl��٠m��*�M�)$GEF��&-���:�A��A;i"��4�W�K"�[� 	Al�Ƽ�/8�=�E٨�GjrI����a�*Z�; hB"�O�QS;����� �?�Q�� �z;�[�=c�L��Y�y�0��Rr��5�����!��N:2��Ce���I�\�4�G0?���#Y�p��Z�S�����6$���?�D�A��@��9`�R�Æ�x��mK��vk�g��{A� M�ټ:T� �M�g(b�]��Rd�C��|����3(63�R񕒛�PM��և�I6L���]y�ɸ@����c��#���	��D�V�3B��[��K���t�t9O^�M���_>��f갼x[O��]���n���w7�[� I��ԟ���g|e \�c����Q0�6�댹�b��ti�"�$J����|���g��j�x
G�l8�i�;+��-�ȯl����@���5�Ol#R���J�xeͬ��,�
��̧��ISY&T[oJ62)�8�K���υ	΋��l�m˯�k�B�E�������g4�#�����W��r%��0����'�e��U��'F�� #�rf���@o����qj��Y��ph�[ȶ�X�Ɲ��B�s亞�0��Lat�B�53j�����8�N��.�������DrN�>ѳ���Ė��j��/�8f=X�^B|��8�,��G]B����!q������U���Y_���3]�Ř�q���G1\W�E�hF&�k)N��6ojc�B��R��9|���޶��T�S�u��f>@GV�Cz&)_8I�a���g6����T�16M��������?p�����0Ĺ],<��I�7[���}�����zl����W{���R1�b�� qm�k|oJ/.�k��������mZ��'����ZL��ұ�d0 �}�>�ͦ7���$�Z(d�P�� &�cHP�r͑� Ki��7��bމN%������;6w 64���pua���Vk=�o�������Lf`�'���`~\A	*��l�{)]{���&��jLT������
WJ����%_�����Z-=��^4��X�@8&^J	��.tN4��62������>Yd����`<YI��}POc�����&X[��cf��q�`
k���	�$JY�D0�Ř��] �N'�}�{��	��c"X��|E��, �CO6}���o���Kkl'@��%߀Z��ڴ�D�F[#\/��v��#%�i*O�Ӗ�����-.��C3T�_��� ��*2���ը��Y[[�16t�9	`	�� P����I����@��m��$z���2�A>f�;��^�˧�L(���J�$e0�xH��4�5u<!��p
���j��:%|�\�)<��sh)t;�����H.��k�7櫾	մG�}�!e8<��=��"�4UuPT�px�O<�)��[�9�PH΀w���N�� �����z�Ϡ�Sםg�v[�3Cݠ�(��O?�.�a�k�bC~�Y��$_!���)|�<��#W��%:�6��d��5n�M�@�z��قA E�	4D�O���!
�|�=�_l��DL���|�� m����Qy�rGL0x���6��%���c���d�V}��Fq:��E�� ���A��u3%��~�$ΗĤ�{j3��s��J�)<y�F:k�f�d�sO�H�}�Ik�m�|�*0�j��MT����N�H���M�IB���@3�A�m��Ld(>A}m���F@����tb��[�l�`��S&��G���J�[h5c��w��TyTa��������~��z���H�qN�� X��	�ھ5هZXڅ�x܉Ibl�Yc��zi���.�J'߂��A0.�����s��DH�����>�f_D�ho+1�Y�r��ѱ����.;ۓ���)3}Vt+Z~��`#���$@�#�W�Q�pQ$H��!�n�d�[/|�̝��Jy�yf��g��
�'�m״���c��fdfp��\�@:���g'��j�f�y�A`��Zr)%N�bB(R�/����.���-�S�,�(����)�(�`=Fw��y��؜i�謂wSLPك�|��ܢ:���)�¥zWw��hA�Ӵc��HL���{.6�
�*�2��f�(;�n_~Yt�[Y�!d��u���N��<+x���)9?)N�%���YVHY�!ua� �T]6�i�1PuZ�U2��;'�+Q�$�U&D�ݤ�I�!�0�k�t�W �*%���(�Н�O��=@���*��ӿ�B�ά��x,�9*���R� �P����"�~��匘��]A��:��Q}��Q� �X b�8ƞ���G��Y���=���c@�>��oMr��!n�i�^L�����f�}t��Ų�p�������Gݷ�&ƓM
D]�S�ڏ������5�h.8�[�����3��D�~BNx)O�[p1t3\LMy�{d-5��gLB�RՎ~��⌜m 4�Ju< �Nd	�V�v^!�NVR\�e�����[���sJ�?�$��5l��i�f���B(y� <�%���;�f�n}3Sy�_V|�؍��tj5ٛY8҆�H�M7�3�SM�I߻J%Gz������.�G@�@�uq	�t$&)|r�����"7�Y�|_���y�@�3�_���.2��e�\�� �I3�J������lB:*�ܮĂ�T��H���u6��N�� 2�|��_倥&��+ �2�G�f�g���ٛ�W2�a�����<g���]c����a���E���$Q�.X\�
�D��Ma��u���1�hO��|T6��7��"2GId��K��n!�����옆dB�v�^4	:�~B=���O�}u��'��;9X V��a��d�cnY��8F�:N��׼z������$D��d=��O��0��=d/Wy�"DDE�
T��&U�\�����&�@;,�����~!�k3�P�؏����\\�<;	-i�ë�o9���jq�������٨����V��]�B�����悐M��}�j��c�9���:�a�{#��D�(�vڂi��^���L�z����������xa $�A���P��J����+����^��/���G���'e8� 򴐴�����n&��S��j�_��lH��mc�����p)PmȽ<p�l�mk��~�z؝T�5���;r��^Y�~�HI�wr&��+#pq������K�.��=xs�)�yA�����;{�i��p��^f��s$@�����n�r������K�i6����>bZu/At8�ʴ�`�aZ;u��R�COv��H�#(4|S�¥��e�bn��O�juг��.��m_�]V+�td��b�ס���0M~��֔�zkBE徵0�h���߸���(�ynO���a�ք�X	�	���"���`�é�Um^dB��^r�]ڨ������E����<К����~ᤃ�����;�Cګ;�U~��b��=������0%�3Y�����~�ğ;Xp�f��KV���-�)�ؐ���qa�|X�<�7�2��N�ʘ��β\f'����]�+_�O��1���/�ef��7��b���Y<J_���فy!j�jQ$�=�/8ɣ b���Z�NY�,>��ͽ�"r-����s��:��z��Fp.�d�0�q�>X"4a�;Lb���^�oFo�0�>������>>��R�����n���'����|���n�J:c��Q���[�*v'2Z� 0���m�,Sm<���^Z��O�[��=]�6S��7��/��d�h<MZ�`ã����7V�*�W,3N�v��,����xa6�!� �-��I�q?��B|�.����3�-J����Ep�L񜢁{B�ɉ�BQd�=3�|a~��z����E֩�������]�\������l<�7����FW��&�����+�̜M�b0�o�hL���Pm�
}�:_��S�&.���� o
n1�.x�޿a�0�{H���٪%���$"�õ��{w�L���<״B#mc%(5��"��Z�d�?+�$� ��s�g�.�dkS�P��i\��ݳ!]Ao!�9���9�c������b����5��Ki���A�b_�ҽ~�CsT�y����2}�A�"ˎ�4�&S��.�OtLr��y��:>�"��|�_`��Q��Ϫ${o/��k�7U�|�������)�8����$>�p`�8zE.G0�;�K�7�|��k�^�#�ʻ8C��Պ~�C.tD����eb��10>e���� j.O2̍!��Y��|�_V�UlAlُ;����f����y�D+��3���/q���b���'��_��4�͇o=�ej�r�f��a���!D?����2��1� ^�Ih��ҁ��y&�UD��裡s��!�-qb�+���n�g�o�D�L����ҏ�6�� ¹�2��c��
iȷB�Ӂ«%�I��[X�����Vs&_�8��K'I�|�ٴ{���>^�Dz^��fjOyG�,�3%o�<�'^}��_m�`4V,�ǜ�j�S��O�\pw4�5�Io� \��%���y|��h2�̓<�В&{�4^L� M��~��!�D�io.XY��ַ]�'��Ø��d����9HE�*�k� $�gS< MbM�HGtwv�Ԣ��_@�8q,<��Lڶ�|�{P���=_�@��)���)��~M�0F-5C��G =�0Y��.;�@qA�y���G�lT@�̶YP��������,��V��=�[�U���=��E�ʏ6�y�=F��P7$����M	Ν��Vv0�-\��dZ��ٺ�Ѻ�d�i�C����s �ۃ��q�\�[���p
��m��ƯLi�wǂX<6D��h����E�2/��T�������K���x[s	�_����o�����-��{��KE9��i�Ø(@9�ZJ��$1M�1.|I���v���eE����X=l�n����vT�����cx.��2�K������)4�IeI���9�+�pr���*�*pV��� ��\�}���L{�)�z�K�|�����`#�2Y��`�#���}���J%Ҥ����o��������6�c�Y��К2-����4�3N��Ʈ�X�G_%��0;e����D����&�V�n�'CRB7$���Ӝ��${�iAI΃�'�ǒ�͘@�d��	�AA�����ul=�(�P3:{*���4t��2(b.�qp��*���W%&���������B�C�7܀1���cr^mf�h}��QS����p���:>n�u���8�\�����X�L`�w��P��wq?K�G�m;�p�p�Q�-�+�w�&�H��T�|�v_��^�Ɵ���mL�E��"�i�a>P�Ꜥ>`[B�_}zt�)X��*#����.��P������ �����X����,�ǰ�{;���]�Әb�j�J=Rdcc&  �"�?K���?�7Ͽ.��/MZ�@�=0�7��y�@ `Fz�-�;�H�r�}���C
�Ɗ�a_UM	��}����@�h��#9�l^�r�]6i�/n��ScCz�� g��4�	��HJ�\�v|�$�O� 1�ȩ~Cj9c�B�)c�7����;��s�'���>��T�z��6o�7{��:�E�����AZ�E��6MCg��IO�d���\<��/��ߧp���m�L��*��ا�Q�7���-��b���wz�9O�Y&N�|��P�8�Ƥ��͋��8%�`��.��ڮc$�Ҳ�v�>	��W�����9n�$21�G�>E�Ԥ	Ϋ/D�>��n	9q3$��1K��:��!�u
��J*;��'�k?лCIO��<S�#�].ƪ�� �+\����(F��B��w�II_��&�6C�� ���q46n�r��;�hˁA��jz.�"%"X�+��Io>ڥ���^M��]M��^=��kPe'K�fù�B�]���x2F1�cT�Pˤ+<�x-�qn��{��[�ǉ�lK�mg������D6+����;3�k]�Ħ�EIJ�8��k}�&�?Y)^�MFL�3�G	 ,}���ܚ�!�U�-M�6��G�2jN�|��;�t�y�-�kc*j��P/�����������y��HrSՒ<)*S�c�)�]�z\�=9����*h;�]���T_�=� F]���T����	�}�7�}�V�^N�t�B�%���-��FO> _��-�g���(���A鉸��q�����]��E���Ŕ�c���Y�4,m����JxN �A�	.��`����ԆI�΋��Ζ�ݢ�&|�}ً�7�k��Oa�Ak��X�	~�!� RC�V~e�[l�:M޳!��E{��%�8tQնPdG�F9�FB�8�����	�c�q$В��L�3j�f���l�w5F�|��96+�uF����{��y<�5c����'p�GW���o���Vr-����D�J�䬱�pl��M��ʼ�㬂MaO�Cq-(������x������CI<K
}����C��[$icaI������Z}�Y�ٳ��G���4�?q5���bV#k�߮�՗�	��w��q�Z�ϖ��d]**��&Kb�����8�>�"�Nʠ�0'�a��z���$:��02��!�6���@S�(5����T�h��TN�	w�W+�c�ڌ�b+ 
�F7{���;����P�@�M<B>���F=���9��^t��i�!����\��g7C4?���ې����%�|��n1Au�g|/y@�m��4�+ӥ����Y��4�p�T�%����I�V�[L�ڝ�=@����J�a ���7��q,�l�<��n~T�پ���d.0q�O\�I=Mk{�x�=bʪ�0��[��Z�SwA����x��gwi�����Ξ _��[��U��X�;H��pO�ZVQ�/�*�)�ޑӘ�n�	�PGn4��"�X
�
�2����V31I'����L����� 5Z��F��1S<�l1���/��޵S�!Є�ٽ��w��'J�����	�y=��r������e�6[��_Q�ww"�Dnx�����������`�'ڸ�!��|:d;o�a��5so5�;�hK1ެ̻�^n�ѕ)%ay�:��S�6���e:��IDo���`�7O���-�J).���z����ej�`����ૐ��g!�q=�clXio����i[�e��~'ֈ��&��vv�G8�+�}�ZH>hj������<L�R��Ĺc�����Z��&gl_��w���G�=�n!ab=�$FVd��|�� ��;V���Gg�{W֖b���,Z�t�	q1e"T�4��F��چ�Kn���u5������zc�X��5��'� <^ص�T~Κ�J��R>Kc*�����-H��,�K��kQ ���O�����u���1��,h�٧-�~s.���������?���2P�
/ލ6P�����،1/n:�zע�XVچ�}ݥf�0�nŻ�KC1XR����mQZ`�D°*�ד-;Z�޿�0���[�1D�Hh�/$M��TCe�L��&��R��ôp�WǍK��R��gǠ��[�����}j�� b��W�}�B{��ݝ�R#�W?P�sGRj,��.oŜ�M/®o؉>.�̋�X�JŊ�}�=�'�n(�|��;e�F_�C�Zo��DĜ�a�Xh$�j;a�#t=�x��$\�}%���|
Z�����*G'B'�B+����c%N#g��ݒg�����+��e_0�L����-+��0�XZs�I+k��m���÷g��k��U�Nn���ֱ�]�C4%7c��<���<���a�%��XV=��)r��APO#��~"*į��']~KN���D��C�����}�1��)�����z_����-�A���X��L�fS� J��i�8c��
h�-��w;�ҩC��$�[ؗ� ��s�e"�|�,'���=��.X�M��<5��5�5�ۘl�4R�@�� c�s��c�"�w�:?Dp�Rn���:y������P#@���{��Xp5"_���'�m�w�u�@X���u�#�䘾í�Zv-�׃�~vU�]�o���0Va��0�V 嶿�#��4Vm@1{�Q%+��z��y,�/R�����)"A[����b��_��������#�\_���TD�٤o�s2VB�<�9��e|
uZ.CŠ�c
'&�0G9�fqp^���|У���?��5 sH���*D�3�"&\�gV��44Y�؊�F�'��_��C�]kw7$z�JHpg��`.��=�,�lsj���̮Mg�j�?훪��ͲbI�õ�穭~o@�}�|pe��	�XgT��q�dF�9@΃ᓹ���d����pB�Q�X��h<�k�IV�s�A�(�k�9ƠQ�?����Z�S�	_)x��5��=Q���	^��*�`�@�t)��e�C��b\Ч�|�p_��Y*^3̿�-�g'�ᅡ1G��OS?�ޞ�����Ią�����W�#�����a�����A���
�'���(2h`w�U!��
W�g�j��v.d����u���E�d���1S0�&NNt<6�ubKd;?��{��ϼ��в�r�/���F�'��H��.�+Z��`��%[��7J��;q�E��
��_F���,�O�.��!bV��!Y���(,Qڷ��x	e�_cK��gS�"�����E�U���7�!��2ు��#���J��7�>9�h�����6�F��s5�����>qML�&Ӻb��r���>��Z�X�M�L��*뷞������yWwCՍ"-3�C96	<B�~x�	-`D0���� �U���_���	��OE y�<�q���@5�
��K=���%�26��Z���o�O1C+�Q��/�n��q��yW�GS�@�X̂/Y�O$���m֎ L�y6i}'���t�SC���*�,~5/KZ�%Xb�-'B�;rhg�0��M�N�Qb'_j��%_���A`������;�������9h��.��0�S@�� ������]�c�v�r�E҆HE�|>F�A�S#��B�H�z����ys��)D@!���=fmL��@YC}�W�����ʅ\�G���I��֣�.[)�>e7�xJ�M�g2�X��1�OfmQ�$���V�q��V����R`�;�i���Ʋtٞ�8Cմ����A	�\�;�4���#��3�ts�|���+�`E��C5���@cE����4��q�l��I��,��<����{��h�	�D��Z���-�q�i9�����/O��/�i���y�����aDGkU����a��]\�t̊۝L�I�_q���oNu��[G��cu����:<�]q�h�|��N��}�w]�ú�&�]���E
;�q=��L7��㑟7�A�* �Xͱt͠%�p�~�jX}����AleCIA�~Wyܑ&�K�Mf�H�ۭ�L����v&�ƭ��m��$-9��"Q��Z���#�j�WAQ�W-��
��^iv�����f�X�L4v�k֧R�����q8<��̊5Q�ƃV6#�^����-�N�v�|O��=4<)����>v�ʰ���Z|����GHe���I@ �%).%l��Mxٖ�P����2��,�D{K�ܱ�$���48CJ��Q(�>f�����p��(��PծnNk��E�J!1A7S=7�%j��.h�X��ZJ�CK�����aMأ�E[�
==��0�3ώ@9�<i
�o�T���0��V���uyI頨s{��(�_m�p�:ړ��4 ���'F����O��t�D�Eg�!��e:�R{"�Q�$l�*�~���3�P�!�E�򾖚�O�����$�E,3U�Qc6J3�yB<���ݿ�ՙ?9���=�}+S
4�bI�A�L%�m�Б���$���τ��)6����Ђ�@$���^;�^�J��1k%���:�'�E(��m*ڌqbg?B'�~��ډ��U��Ӛʓ��;�Q�`��{�	��<����9	�O�d[*�)�a	V+�%��px����	�g7�z��^�Yo42�%8�A��w� ��N��%m���!�p�����b�<)��N�~��Y\rQCE&�S_ E��i�x��Q�Q���i�}u��!�sL��[��7���-`�' �I#�� ��` ~US �ah���:�ؓ�o������h�-&��~'��Ѕ�$�r)�×?�h�a����4V�Uę�~-��%��2̗�âc��<� 6�c�ǻ�j�M;�����<���ny����{��rl-֎���iʛ+���s�	�:�mkկ������>,Xuh����̥�%n��i�r�KR��V����0�պ�ֽ�*��!-���c
�L��޻�t�?-0R,-�ۅ�s&�2�"b�Jy�^��ڧ[F�b� ������b���Y�:l�!�ȓ��?�a.j�� �N٭|�T.�r�����IH^�];�6b�V����#&�\)@H��j�2	]�}N3������	�l{\}�BS������ʮ�� N���Z�L�����m썚���@���j�b�\�b �$ׅ���a�"��g$�P�v�z�]���`��޼��0w235>@`�����y.��t�u�f�I2� �%L<��2���o �����m�_�O�Cu��"�js�	1��?�ͬf�*I�x��%����I��HӽS=��2��Ѡ���� `+*���1�(�L�uj1�u�Q�g�ֈ%��:q�܊�~ ���XF��_�"��k��z�kD���C+-���;��_SU~��o�A� �x���<WcqxXﯙ2��#>o�`ɋ_$�ץ`2-Ɣy��8;2˥/���_0(m�nUL��\�=���AӲ �f:��O�51����A�
�\���~��y������MtO;��'o�9ULv�k��1ǃ���ۨ�H�b�5�dЛ�w�D��LeN��K�ѱ3��v�(4��I�W0���c��`�V���hP�74d��m�/B���L�\9]�͟%�$�=�����.��|h�����!��侚���
8����]]�? ���͍������r���6�4���s���菤��s�E�!j�s�e�Ļ��KP�Uv����y��GC�(FZ$��y���'A��
N��,w�Tq����Z1~�����`�281�0���
��1/ɉ$��^�0c��0aO�*���ޘ#8���2ʗ�0^��N�e�,"$�UR�yG{j�6�H~J�՘�	����OWt6-���lL�
���J��9q�/��c��Ŗ0��,��(�`�̙0z{)
�+JU�@�9�_P]��Ĵ�T�<�����r���@(�JT!�#����I����f����1��䃢��Ɓ	���:������r�{������1	q'��(r��cO�7X���b�����j��b���g�B*�%[����o3���:]�Z&I���mi��cس��*���x ��ck���P�C"�ܢ��8����if���L4>�@a�s�v��2DSw�>R##Ix�p�z��$Y�I�^tf�.�I��+�9� X:I�}�D�S �� ջȭ�¶b~�,���&��W*��R4�_k*$��������֤UD�QBRA>ڞy��"�˫��My��E����t9���m;�Չ�B����?`P-�c��P�;��}�ܪ� �}��O��6���i�Q�r�2��YgC��� �)�_n��e� �yI~�i��;�\�,�_��
]a��N)�5��RN9Hb>B��m���)6���+"��ge�����o��@��̮�\�~Z8�����_��a��~P��t�}7X����N��	��H�T��gH؛�c�����z��M�h��=z��Myh����Fx���t�=k�s�$�R�q^��V����}�7E%N�*�����2h��3�ڽ~4jX{�qo��<Ýk�S94~#͓'X0����䥝,]|#����(��*q�qk\~u����o��*/�l
���\ ��ZbgΒ,]���]��;\G�?��,��}��:�!��Ί����J�%�Έ�,�1e3��+b�|$��4kt��0��c�4�NV����⦦蔃��l�$���'f��F�&�����8 �*lo�����w��lԋ�3��}]:�:�v���6�ޤ�t	�fɗV��l���f��[���?@�hk$�U��>����&އX5{82��j��^ǧ@ݩ~��ipe�\I�zf��j�o\�E��!�j�r�'�u�1�oE4Wd�m��38k^22�P����#ְuh����sY��b�aW�˩�.��]h'1�%�A��Z�R��'`ZP?�>�e�c����Z4��FR�ׇ8#��n;E��ے����d�P\��S��=i��7\�r_y*�4(�4��V�9?���tQ��>!�f9j�,]xK��D�E>�m	�Dz���T�i93�8�7?���z����Ҙ�t��5B�3��"!�|�G��h��I���Xzi��	�2�9��Q���'P��!t��օ�����8�����G�^�/�|��Dɷދ0�9zw�d� �O��j�?�E�>�7�}/I��m��u�4Mk����h��7-\�w��
7$b~V.� q��O�z��'U�c�����k�z�������������'s)6-7���7����cV�3�)�c���|Ao��)'���wh�l���C7�e9�hQ$^��M0��l�x8�A/�j��R���d�T�F��������.��Y�>�c�Z�LG��4V��N�0܋�l�	Ry)/�&h�w��+�[�ojbn��jWv�N�b��QVE�y�kA�p�)����6��'""�hi�\�F�TZ��PaWs��[�2�����T�E~��i��OB�~a����¯.0 ��LΉ�V#�em2-���
B��u]����`��iZ;T��emo&M����t}��Ge"͡&���wH��k��x�b:��)��h��P@����7b��w��P(
6_���g�5/d�`7�5<��!<��5�\k�x���*@z���6Y��4Ԅ;�?>�/3E�BQ,���A�
7��9'_(�$K���T�L�=�N��a'2���iM���1��X��$@vw@b�@�U9���xh1hB��Z�m��bh�5�|�1��%��d���8��!c&�U�H�OL9�A����w�h��w� ��j�,"������b^���~ڰ�LvZ/>OcSn]�e�2us�v��i���7{3by���*��a�����*��t�ow��G�,��~jWSi�o��u���b���ϸ����윧�v`��"z��SF�ԃ/�&��S�78Y�t��ε�oM۶g�s��=�@�eާ�i2�L�'%�`�uᩳ�Bi:��I&�	5�Oᓤ#EiJ����*��ex^�׫�yϛ�Ӭ��ᨹ��V�Jo����0o�_N���#lh<9�qa��a���'"����(��)�ل �9�5|���A�GEAa�O��P
m�Ƅ�,L���S{�D��[6Uw��ȗF�=�*LU�g�����I���?$qv�s����e�J�Bbj'�z�ߚ?��! �9��_X��-���P�U˚�R��o����F��oq���GÖɝǎ-oI��j�%� ����^�f��L��1��}����� ��5��6V�!�@�B�f�f�Ko��ES�y&��`�ap����w* �wx�C�6܊��ke�f��D�y�QtS�`��,ʖv����[��X���ڦp��'y��Q�Y�R���.*�F�_HCA�=@BZ��݇�D�����C������k����&�ʲ�sv�a�7��\cq��PV��cjY�=�>�o�8*����u�vl֟۸ĩ�I�3������Rmg'm����*b�>�zMd��k�]���]��5H3��1&\�$q!�ݔH74�ct�/:R�3��E�P�fȊ��u�T�.�_�}z��pz��h1����>n�!�" �f̖� �&l�r����E�ا���)M�L�ȉ�F�o�Onq�򊅳�Ss dx�#���U�}�Ξ��EMb�g�K�AC��F�����r5���h�?��īrf�a���Yz����K:(�ק�|�>���!}q����b+?��6�!�=`�P�:g��d$�����%�_̻���"!vwj�(����X���,�+v��>��IZ�N�p%�i2;�~�kr��{�[���kNSY�-R�qD��l��Ԝ^�@{H�𮔩S��I]��1iV�K)F�BS���;|�T��������x+��" Gq���"m�o��
J�|�9��)���6}���EZ,=Z�ɞ��V�/�3tiL"�n�=nF�
�}���a��9rtq*�� `��w�9��}����W��jxb��B�e�eJ�G�!��,(:-��k&�{FMag�A�,�?�kޏ���$a">�3����l���	7��g��T�^n
@M|Z�<L��18��}5��B��F�IX��fBz6�xd�k������/��'5fo���~	ݨg$V����?!��RO��m� ?��y�(շ��N�o�g�)vc��v%� ���e0�K����ԖK�دN�q�=)^��+sS�\��-�Z\���i��J�I�a���6l�8󫳐��#kII�}7�?�A��n��Ǭ���:�T�V���<�)Y��;��n+
x��qܹˠ~|���L�h*�W]�I�J�o! ��a��c�n���Bl�~/��K�˺
!���r��������c�d
��kpW5<z&����/����^�'r G^��L7ϴp`%3$M"S��"���xC_z+�,N�UYu���#�E�Vs�.��*�y��'���Η�qr(hW���4�pa�����w� �\j �0b��� ����d�&�-�`�!*�IH����jݮ�[6���hUT橀Z��CU-	QD}���	om�c�WE�~�RG��^���>�/c�k���2���V7��1讃̳eEm~�3rq�v���}�%B�z��>K^�h`g�5���M�ܯ�����Y��>���H�80��6:�2Fdu��nn]�Yl��Fl���s<�lzk�L�Ms�Y�J60~�3<],�͒�A��kwym���A�V���hj�U�	����l�����#�4�G��-<A)�WZ���CQ�����>O��p�{��7s��R��'���](����Bd0�}�뫞�곀�+�p�����R�9���ʀ�])?�f�D
r�y� �GL&-"�j
nMf�BMM1}�&�K���3>��d'�b�D)��ǟ
�oa�Ə�Ij�g��,�\��{l.��]�^�[�صҕ��;��R����-s虞��V~=�Fp��}_ˎ�+�K��3�$R�ă�n�/�~�!��bLf𲳇�H�ws���e���e?�W��}z��Oy�LLču]��.�{�I�|F�)	����8GP6ۭ ^�g���jCI`L���m��4���V'Q�%��\vضU�ؾ�W:����h,�݆�/�"k2���gL���ت�9T0�E�����O�Y>~�$�g���d��z1�H�K��=ݐ�RR�g'�L8�8�
]B��Y��x��b̂�BZ_�������A�W���mP��!�P���ռ(c���8H�����^�k�ƉM���m�'Y�A],�k�W8l*������Н ��1 l��3'�J���c�7���|�`d���u������ �;�Ҡ�T�ba��M����`�cix� fЂj�y��%�t�X�R�`�BeZ��Ѿ���]�o�2���BI�7��v�"F��vU�S���J>�@k��-`���*!Z�ػ�}�'�/�pv�v70ߛ�=|��#��C�����R����Jݷ��j-:^5�G^��O}�H���Ⱥ'ȢKe:����n Ia9���o�g���F
��8dk6N� w�3j��5�[�_G��X4k��"Bn(~bnKh͓GӅ�'bT�{� �R���|��e��I�N�쟯O�K�AW'EaQ�;J��m�0�۞��� 8�n��d��-�WF'��[T��g	���D��K����'g��ǝi;+5�sf/�
ʼpЂ�t�T�։-��Z/~<���i.���/�v��N�K=,����cR���t�G�;����ld$��B(���9�[�:(*^�U�����qn����U�t�a���(᳡��<�a�Qy���9��+�hܐ���=C��{+F�(��wі	Y�ߪj��%�Izd��L�.�Ȫ���:w��@bIg��k<s��5���=R.�FC�~>�w[URe0���c,�� �@)I�A�w�J7Dͅ�ϵG]�����aި��R���U+�7�>'��+��}ǒP�i�18�o(�v$�8�Ò ~+f�u=iD ���R�s������S$�������,�Y��G� -�����h����?{3�=�b�`9\��J,>H?4U ���?3�+^7��PGN �{\�`��C�HO;��j���wj`��Ǿ1rf���Գ���?���,ڞv�J�͙D�Z~�c�$�Xf�8�^���qyB���C�/u��em$�QA�rV
�w�/YΈ+MG[d/�k��vsOF���Mc2F�3��jL+.�Z��>B�����k��V3�1�J�R8�*4ȗG�e��L:5�/�%#|���,<^�8����.C�w����]�ݝ��`2�`8�3Ѿ��Efi���}�y���-F��m�'l�,����<���`�S��@��4��|ػ�t��kbW��bF2�U1Ìm�]�������"��Z�a�u��R��x�0Jte����!и�I#�r��_�t�;�/Q�帐-s�:����#v(d�Snr��M��
�Al�9np�^Q�@s`��CKuC?e�2�����#3�͌G������Ge��͸�Bt`�.�Y��M���d]��� S8F���Ħ$K���Mſ@��k�ē������*���P�+l�!��]򑆅8�WP$DqxBf�:�7� ��5��Yz�=:����&Q*Z���=ߥ{'vw>�.�jM�4`�@�d��ǲSԓ�n��j�;�b<m�d�.�lS��p/⌸���,�(�x���
�����G��c;��O����?q�y���XQ��|A�)�q����s~�+D7O�%"�Y%֍c8�u'�Pzl��'Jc>G�֘?�^Ua��%�yP�ͳj�W�FsLo��F�y�(l��Fj�
pկ��+�P"h�x*8���K��ש�Cǹ�<�Oz�r0.�;s���um�U���֜�ǜTfB��Vv������ߦX���FK��<ɡ��צ�_ϕxW��6�������[�039'z�Tf��s����Tr4G����/D+�~�|&B����T:i�m�DvE��Ōn�W�zL�i#c��\�w�=8��F���o�*�+r6 ��KL�)�k�a�����k�]���+��.�
Ⱥ>nEa,�ꭰ�:G�~5�Yocx���v��/ ѝ���C���׌�Q�%�+WC��j*Uހ�	���E)!�A���׏i���J!?P1������;���ѿ��"�5�,-[������������t{q������\3\�I�q�1�-Sp$\���v<�N�x���}.Z���ƥ��Xǵ�� �x�`";7T�V��ж�ڊ󤝪��LӼ�伈-�޾v"��!j��{���<-ۗ�&��و�+˶��a��z����mC��̵�Wt"�V_k�d���G[��L���b�\���^E�Ų�~����_¿�7���p�˶�y�B���#_IӢ�q�*����5�9!���W�sw=��q
z)'&��-7Sbci�+���}�c4{40�N<V�̨n��k1��B-�y�ڑ��(�WE��Wl��=�fO��l�6�=��Aj�^�Z�9ug$������Kn�F5��.���"��婄@' �6��7�n@�c}�ǟ��y�h�ÊA.V+����+�1��j�(� ���u�������N�~�/��I��!WaD}���6�y�)Y;�^�Cv�dx�qc�g$�:�bi��PE���R ���MoEsTu���p�N<��b�s�C���吼hf����[��`֢�Ki�'��O�aZÖ�Ӵ�Z��K	D����j^�1��d��0-��i�ݝob��h ���,<c�O@�*V�̟6Q
�9y��-�`��|���x''l]�C_�߻�4��ʋp��w��1��-��U��hw���ӵ�+�e��9uA��K�wö�h��~�FVC����X���`��I4����P �ZD��'"�d\V�ps,l./�l���\���
g�dy-'��c�3�]���q[��[ߡn;�#0-{�_�GN:�pH��Y��E���=~N4~�O��R�;��9)p��	���W�W�
c(���e=����/�SEb}C,�y�7?-.��z���ð)m���{�I���<G`"Ǖ��i�6�-�Y�m��UU�p25���F��A�f�����&���{�|���lu�
/�{,UT�=�𵇔�r��S����e�ve_I�|�Ve����9ʻ��ƽ�>�d��%Sc���w����h����g*k���� �S('��� xF�|������?na,z2J{�sD���6:w�vZ�5��+y��E���"�s���C�Gr��@�9>&FaQc���bs��tK}Qf�\����i���DV��[&��;0K⫷՘�fre��$mq�JVa^���O9���L�0�RXr��=�{"�Uk	ǽx���(r-��n{q�$�=����7�Z=~$���>ۿ�$��>������`if<*���0I<�Ľ#����NRwG�޲�sp���H/F��@h�6k!ߵ����,�d���;�2�����^>�"���yC�1�}h<@����	տ�U�Y����F�Ӹ�B.�j���&�?�����ӈ�9K�n�衇1��Z.{�g[������܊�̉}
5/K��DN�3@iwx5���#|��v$62�4�L[�Kɐ�1/���{�BR�
1��y�v!�ABsl��P�z��B:T���K�XQ�#i�A9F�l�oHbkD�w�s��͆F��6��]�h��_����#n:�ַĜZ�� 6�!yJT4  �>�{dUn��o%٣�(<����J���މsn�M�~�k�u�/F�����{��V���X�3�D&�r*�#�-q����bؒ���
�i�>�߲�p5�@�H�@��P����tl��=H�Հe�(s�_D����i5>���ϴ�/B��0�)y�F"T�ܪJ7�Z�����7
�_9	<�)RM��X7�W@����Y�]�J����	��������^�,�T,"˼���L�J0�7�M�\�f���?y"�|}(���f� N��{�r��Q`@��}��(P��"hCݿ��w<߆��M�;�L�+�;}���(2����dN�{�-��@Fjg����Ě�Eꖊ�',;��V2ZiT�i=`���A�]����:b�aN+� u`�������V+vs�mc����
fSdv�e[������s}[1Uҏ,')�8 �X=�O`���dE��-�d�ِ��,oiځ��=�d�??ڟR'��.g�?��+����("����	�}���������	X��#U�7y򮷿SG`�˫���]<�X����ډRw.���&k��7	�r�lN ��B�IB������K��#���M��[��Xtҝ{J��=o�����x$����(�%�'^�F�zQ�ŴK���aU�&�e��0���V���Ȅ��C���o���w�GB�:i)�`e��F?��a~�f���'�кkN��h����8rn��y7���өhuy�ix�F��v}Q�ԮC���թ(e��n=��H����B%�;MV��F7]K�<��e���&�hM��Y�>?���źg�k��4Z)�U9�[)�gn<lO�@�7,*�8d��}g�"�)��0����J՜}��mf��Z-���Jg�sD2�H6.�0ɯ�� ��zdk��p�v���[��_��z HJqI�S�f���DVwsS���T^���(wW�k�j��Fi�����G8��W��\L�
��������{�s:h���%H�q��;�{�?v�x8cCm�/�D��?�9;��+	�J|�KB���՘}�!��_��n#�GZ�$^]©���o�G�t�M?�غu�Y'���:WJ�&F�)���F��d[3�5E�ht��dB��|�rr�tV��+٭Ѕ�Ȉ��#�v��!6�B=3�<O��4�'��I�����zw����t4�om<<K ��X��&g�o3���Mk�������~l�xZ.�$�I^��3^��Q8����a�>$wa����`���HT(] #ZV�@�]੣H }Ҁu��V��V�-}x,���=��gw�@��ndF��F �*��J>�1��)H����an
 �9�j%Z�Ɂ��ߴG���?Ǻ��e��"�x<��l�qD�Y���.�,My�O�狻w��8H��}kzf:�j8-���/˽�<ާ��ңˀ�<���$"�4@��R�{wX�|��
a�|Nq�i�k��Ӫ�)цL]S^��c$|��4gM�(�g�~�_���X���9�?�t���<��˗V	����Q��ʹU����|y�5FBRs_�J/ʚ꼒�$�(�
�\�g7�q��v
�*&D����-'9$�X���,�	�<�3ƌ�z D�b�#�t��*�$�1)D���K����wӾ{W2j����z�b�a5=ah�=9�m)EtlBu���ص���wቑV8א|��WŰ�h�jc���)�B2��F��{g���4��3?'�a��u3%�	~Q�qĹ���Փu���i����V	2�M��l,.K���;��ُ��z�5z�����z"D����b�l[}�4�a��m����"W�5w��OG��tQF�~L9nZ�,� ��Ͱ�{��L�E�W6M3Pi�&P|�kwF6O�d4���1�k���l�?5i�I�՘�����I���rf0dyǀ��<'���Q)��2>A�*va�QN�$[�,�������0�;6%�Z�Y�����w�h��S����~����xX,�Z�h����B!�s�rK�m��oT������1��<�����Y�_O 分%���� ��;�a�5�vA�iR�~�{��ĩ�Kt.�ݮq�V���1U#L��~���D�%����~Ћgf�$�R�t����tx05_V���Tp��������^b��稟�s�7�������0�Ԕ�Ɂ[^=ML�:�	����g�8ɹ�{���
��&̓L�kZ�������% b$ye0��>A��̢[3���ӵd��eB�~�-n�CV;�>o�i��U����]����ǆ$�f$��ݡUU����r!(�]}PW&4(�^�u���~�P����e���~+��w���M��۰&3KM�N�#�K�~�2N�MH��ݔ-�Z�Ƶ�:Y2��U>Z�x��W6�'�}��*̫�l��=�O���9��ښ4���B�-b���B?|�B$���R�S���z�4Kĥx(����ޞ��)�ѽ3�kQ=E�6��E�"S�b{�H�mx*9�(>:/ڲo˿c3ג�:��T���jj-kd*q�##�7>�����c�Z���Cس���J����gxkjl�W�~jY7<�`}�hvԗ���Q%?[��?��vN�ח���&a����p�s�j�����t�S��:���:�\"���̐�|�E���A���=eQݵ5r'�e�|�*�~���v��x�'�S��^-��*�J�9��.ҋt,.��>V_l�ьz$�jV����^AJrT���,,�L�]��pI}`�B���:ˤ���܆a?���is��9U�k
��1�KZ��s��wI�U���m�b�	 �t��N���3_�����e��zZ�SrA���Ԏ��������[ ��@�ɅF,������Fs�|���Ѡ��r\�l�/�>�����k��y�c��U|X��im�9d�ߚ��[���/g�V�6�Δ�'*#��WݣB�����>�I.d7�95�d��e������6��ۘa���.�~�)��^��L� /��G�׊g�;�>׋�Se���:Jf����5M�������Ƚ�'j��8p��p�~hl_�2�ŪZ�C�!B��RC�e����+�**:uL*l;�wLv.Ȱ��c����~��@Uuz"�
\'u*��LZT�F�]�$�TZg�P@x�JE}�E�c�.��@��?5vlJ�����>	���55k�o(S������2��rĕ�}-��B��+�[G�����;����0�MO��v�E��yOJ@�9��x]�%��w�C���E}�S������h���?�)�fP��$"�>g�k� ���/���`��<�uyԄ��F�
��Ek���@�R(U��7O>�P�I��NQL���Z�����L�<j���N�X��G�}3�XM(��5�YD�t�s��x)%�(h�����>|���)�G(s_�~>�e�!�$첅��F����ńKX���M���p��a���='7
dw�M��Z�5pn�_Uָc��ao�*^�Ӗ�b���k6��7ù�M:��]�w�G�z�Y�\�	�~��?����x�-���1�8�q�!~Z1l����I�nK���)#po�O}ZL2����?�vF���t��5�������O�x]J�Ən�#ED��#�&6����d:f���GTgջ�Jm�g����@�x0Y���E����%s����l#�UE����MxE�n��ݏ�йT;̮3��bYŌ�`E�Kk0�l��C�U@����7~P�o�aT�5��nB�;�j�O���7�Z�u�¿2*��/�4�������'��NT��0��iϹ밍C(ȿ�,9���	#:P�<���Ds��(�}�R���Рw"�6��>�41��C.+_���p��T\�˙䅪���I�5ǕQ%AO���Q��*�X�_�"*&�"V�G�x����V����s��1ԩ��,'�<��&Y�J��N�b��>��W��b�X`��BBaP�G�Q���kkt�l���tl�uzV���G�$Oo#�)�ю�γo�m0�����Y�V͢4`	�ⰴ���1�s��_,�rgwlOBk|2>}����v�tv�R��K�>*4!����ܔ[x��J1k;�4�Q\�1��N�����g=*�| ��h�'�N�q
������dݕp뤥�����@w�̼0E6��a�l	$,G֢S餐� o&����yj���F[.4p{X�E��`EAW�JN��j�&�YGЧ�}9��ijv@�B�S��v�Z���Q��I��c�g*!k��$w%�_��sU3=���YKڸ����{�[�aڷ�+d��������O�mM��w����[��ǃ�	!����>R�>����c:����6��?�cGH�����'r�� ��E`7�\E�0�nA��w'�k%�-��)�-՗���3�$��\;ձ3����ටp�.�"�/���4z��*5��9�& TI�4��=@�5r���F<�Hܛ�QJWo�X�ʙ�a������a8�[:H�+t̮����"�Yޚ�����[aÌ�2�oMWi�;"�>��da�<^����Ղ�1��ge������s>�﬿���^��F��D��:�6{˜t^�.���Rpe<��Ġ���8;��B6���"�R>�?b�3�G'�̥�m����s�pdk��Uq�,�9�;V}��ha�$θ���W��c��ݳ;�p���Rs�TS�X!F�o�ʂ\����>g�o�/�]��D��[s&%/ţ��^K�Dq]Wn�5�a J��M`
o끚�1TeoϨ$g$�?FA�ԋE� p�c>x�<�̀�/vv��ˉL�C�H��A��	#.\p ���R��Ȫd��j�ݔg)s:pÊ�0L �.W�LH�x�
���]n�؀>�FH{|&��fjq�J��^!����:�
���a$�Q�'���g���	�ʸ0w���$�����/�{#~ao�?�d+�E��Z�A��^�f��Ӳһ�h�n���6����x����&�I�D!0���}�gO���Q~+��}�Õ��+� �R`�y��|��?VY#a�}�7����BA���i#��0��!P�f8&����'�*���Z!�m ����p"e��e�[,eE�{؋�?
�Y��g������g���$D�9�Y�b��2tm���ީI�t$���p��9'ɻA[}�������:�Ö/o>3iURs�"AV�=\�C7�p�D��b��K�.d�_�6u� ����#���U9h�,3xt1}���MRf��-M�����.��ت ���a�vW�������P0�����m��3�>w/HE>N�g�}��b1�]�R��X�w`��T����,ᯁ�2�;�oεI�C�)P�t�{�Ax��sA�����T��*h������>�V����1��']w,�ye&å�H:kJ���Twb���W�3nv-��r���T%�q���3���%s}c�����.s�2-��O�QLT�1�D��gs�T���P�.�X8Ff��b(�5K�*u�#��G�{_�T<�$�rl�=���z�|"G_��G�g���G������5�<K�|�a	�b�@��;���.�p�Vo��� � ��m ���#ZZ+e��ߌ���"�� SC�PUr���
,���������=�Y0H�������Ad�����a.t�����`6�DP�&�P��S�5#��o�%�V�p��7�"dŪܠz%���A�'�8k⍫�����Λh���$Lep�x���䓊M��"�d�Rhd���t�*��t�o?6 :�|�B��
i�'5:����>��B����;�2SJ(��ݡ{��co��9]�+7.��`��S����"p�_d�J����Ճjg6�U>\�1�B�)F�O�&~p���a�!ky���σh���0껥h �a]o����[,��K�v5�a�҈ �8$<�'`ߋ��z͍��b��Ǫ�5��H]�ty���1*����|e�{>��R<�l�:�q�����k�:��(\6���v�=�=߾�ܒU���a�`덒���7����_ǚK�B�X��,�+��g���7{��&�^&�%&Ҏ�br� BWI�Y���@��dŬl��J���̡����l*W����+�c�R�}�:�Qstp�H�nD��>S����Ca�sl����=�f����wF7�v�u�~�WIR>�H0fvL*�y�wЈ�$I�y+-��0�ߜ9���>Xm��خ��`�dKRY�(�ʳ�>��U�Z�����8�.p<�$��W=�MW������"�����sW#��29I����c���ģ��S���a���۪3���˄&،r�0K��d�^��X��y�0/<�a �_%`��e~P��@7���g�D�o�ZQ>�>�6PQ"]�ʊ�[�PA��8�t#0�?;U���o�k1���qm!>���z���.)b#�A�/�"��;���ڛ���Ä9+��ޮ���#�#�I�c�e��e�-���k�-BӜ���\�*f�k8�Y��C�p�1���0-z����[8���2d����+;%��**�d�*=��r�I�@����]]����Q��r򘡜�������W�cy�2�⋂C�;�恢�,��ݭ�v���N�y򃠏`�U�y/�;E�݄U|�!J���1��HX��=���;�D�h��1��sTv�;��w@�3W�><���P >QH�Vm���"kho�Ei��bK��&���f��Zૈ�H�$MH���D�������$R/�1q���Մ5{�p�
=;�*B�N�~rMn�I$��c�\WHr?���l1C�N.n��p����@M�	GQ�g�e�
X\����B���(�����&���Lƛ��RN��<K����Z�қ�ϲ`�9�JBǈ�x5�]�+ ���Ú�_/(qgԗj�9|��9��:�Ԉ�?������d`��}���X��"� ��d�s��Y��y�)���m��.��ۛ�0��s��YV����Ę��{�{�a�UX2M�q8�zh:���/�ҝ��7��q��I�	�%�I��*:@Ӓ���E堾/ο�b���a�!�diG�`����V��2���DJ�zZ�㔂�Q#�njN����ⓤB ;����i��@�qϫ����Y�{�a�Ɋ���8����f��X��t�i���ב��.�]�1Q��ٚ�I�����X�?M�w%s��}�?ܒ��==�p2�qh5�x���t���W�/;��:ja(�U�;�'Jb/�=P���"�Q�w�����<��[_#M<����[cY,��D <؁�@��p�0��Ŕ	` R\t����Q}w½r����S!C C�Z�	��RX�B%I���
��<u�<�|���\�j`��KuK�$������A��HAI�ꐂ�*@�
���E�x�ӱD4!�`PV��\df�}����F D������R��V���v>��eZ���)�X�y�+�`_nN��H�L��~es�2!B�!x�~��M%�����h�Ծ0��G�-��J �Փ�֘��&8�;�$"P��B�!�yi�/���w�t�á��io��dpڧŒ��n~���6	- ϰ<\�u���������܄w���y
�ϣH�q���;�>��Dc�~��/����n~v�����!Ug�}-t3>� �!w��q���^Yk�F~c����쌐�����Iε��QQ�5���"��|g��b������8H���b��u��*��(A!����.��x����Wr Ͳ�>wY+��2�5s�G��[	�qwvl��/h�	U�x�َ̭̪c��UZju
�n�1� m���O֭�~<��3��t���;��3�Y�����a@
9�H��*(z�=�CZ��?�[�>� *Χ�L��@������?�������w�YC�mR� ��'lU&
���A R�X��c�DK�ڰ��;80�;�Kͻ�,�)sw�7�,ll� j�#��k��Pg>���1�`
����N�6�i�� c�k�	Ri��	�0��{����>o�ǡus��M(-��;׃�0�c^�9��/��R��W�5!�uP���<~sS���� �����}�݌|��_����Κ�̥A�J^�������s�J<RSҍR%�Z�b~<q�|tg�;cj��r�~�k�,��Q��fWt���Ifc�A����H[���Lc'�n#��c]��J�_��N���푵[�u����y�~N���^�68{E�	(Qs}���������Y6�[R��ʊ^���#3a˘������2]�2'X���7',?�"�v���3�kbq�g`j���*:U�S9�� Y��sXb	u�(|2�O�HE~��q%�N�I�$����i��97��'7?NX� �C������p"|�=����I4[�d��+<���KGppq`�MA��|�G��>����£��������+�b�u�ڥ��æ�����Ag������WDi^N�����}m�h-�欅�Sl�z���S�L�n~e����G��]��N�lT��N�^j0��O1�m.�F��oV�Ľ��WdZ���n%���o�T;6��ԥMa��v�P�.%TyB��U/. ,�<K�����<	.�,�\#�֖Ր�:��Oh�w�-~W$99s�S�F?�Q��k3�L�0�/���)���k�nW,�m�y��x����!8�a�c*^�c�/%pk]ަ������?��3��Z\R�J�
N��'	<s���C�"��!��!�3���I�(_��R�|��%��˕�� ���0P�L�z�^�_�|�P�#g���}voS�2��xh��s=b
ߍſ�u�0b�'Y�Q�R	D��y!�&X�U$�3`},Jl� ��3�jFgs#c����¸����nLCS.
6�q�k<���q��$��pӆ���/m:1�T@�N��(Q� Q�*<z-=���&�E�T���e���T�.�\���E3�p%2c����K[gk���z���|�������vȾkN�$A�l�â��x�FP�(),	_�K��_&�1L�N5jس��4�$jaj���=}b��h(�_h@	m��Qp@�V	��/�X�e�����39E�J�B_�B0r-o x�B�8oq��Q��[��=ڨ�e�j}�Ǣy]q�������q�`�}����zoY�II5a���]
p�!�[/��+l��!(E�=��[&J������+�ʲˀ~�r�qn_���sa@|��T|���9�KSm�R�)�߾�0#��bF��]1�YUk y�o,6R���?g� ���Zϡx�fEgP�s.\J��N9�&�����Z��1�]�^��e���u��y��alx�hަ��`ј�!ߨ��<��	��(V�}��\<i�~q3��y��~XHW�#�ZU��(�Z�d������b�6�o�x��}H�P�`�w����mf�z��-�O�tIq����/lq�2�e=Q�e��.>	i��P(�pC�GQ4�w`k���+|H�����p�x�����6��W�
<��جl���}����$Hy�o��=�bi|�1��Ut$�6�Ѿ�9�E�52�
p7���.$�s�%d���ʤ�.y��{�"U�kI�iݜ��S|���F@�,����gO��j$��6Ӊm�;,��8|�ɿӥ`�1��S�\�DX�����%�rU������C�rS�
�B�a�^����HH#t��lzx�5���ŗ���p�G��e�0�� ���ٕhA3uQݎ<yt-�T�;G7�i�����)0�{�>iI=0�����\�t`*Y8���]Pp��U�ĂݞR�U5E��\��\T�<�?ů��by�4���1/�����Ӂ�ghV	��F]"�%Yl��:�w.�T�>sR��g��=��>�<�ɘ�V:mo�J�7��������V��>ɚ���)_��bIˮ7�F�V�s�X)i^�%���4�ڂ�m���KO��o�Wc�ہ"p#�_�_v��!u&��\�Ā�{�Y�p���kB`R�&
<`�?/O�����,Z͹���?���uD�飬I=��P'�� u��$�j����o Zb�lؒ�ƥ\���$������E�I��[���$��j��Dp��iy��B�8P�)�6��1��CC�lq~��p~�(��W��MD%?�������I`��4aW�O����Г�j�a��hl38ɺ�bXJ��E)<[P��GS������?�	� ��o�*�����?=d�'��ܖϰ��j$m��@'׈4v�ǚ��0�OYJ!C�I�+gN�g�3�&!/[��>	P|lv��$�)���Se�(Q�Υ�ڢ��t't؞�伐>���W�f�����<�pkte��2Ԓk��U�5�!��|�5��H9�tN=/�/�V����K-� ��B� p�X��"f�×Q,�j�E�}������(f2�}M�{���>�M�*)�[Y��#������1�(���s�������,y[��P
m-���o�+G��h;�{����Y��<a%m��!8�ڷm������	`���<^�b�v��(�6�1�|�g`vG����QH3�H5�=<
�3F	<>䎛�a���w%����4/�㬨�S/]lc��8�T�-j3�����pDL�<�łƪ�¼�;�1oybP	܏��_k?@�rk����>ز_1>����	���O[_�V���R d0Oi���A�z ȝ�$�
~W�=Q����kQF�ٗ�Z�K3
ùʽ7���sӋ�K(�5�"-b���Z��o�E)�s�� ���C�.�c�%�V�i�Ƭ���q��;����+���t�ި����9��lS�5�TchŰ��=,r�x�.�T�%I��	 +�
�,�'����Q�E?���8_u.i�Þ�=��ZO"*v^d:Ԛ#ᵨ{_��r�*H�����?X�ؽu���ЉN���~���݈�[G�L`w�k4M�m_�D>"�Y�~`�.�3��]i2O�}��'���Vz)�$�a��E��9v��=��@�+;L��΅@��'���ȠN��.��{Ln��8f����
�-���|�(�����(���R��3b�KϞ�	L<�����fYK�W<�;{x4ݵ���-�Wh5#��GM�O]c$c8Pbh�Vݺ��49�;&��e�C��Q�����/�-;�ωZTߦ)^�P
�z�M�XO�Y�|��XoZ=�=��<>}��ԙjd�i"�y����f�A�w����Yk������m����h\�K.�2\NC�7���GT\��Pa&i�����m�x8$��O})�n��K8�]�Cxg����� r�4w�dJi֎!�l)���/��.�4��n��I��P��07�eg)m�0�El�8���Y�C����L��� Px�H	����XD�D$�'��g5@
y*7�u������0o;T�U(#���˼��A�ޡ8t��;�r�����9���.:����Z��:���	͉�\⁷�ņ�����u�$�Ȏ=�
.bv�)��$��Du�z����AyN��*I��\r���k���/9Ѻ]A�����\. �Ő08t�)�:"����n?5[�e,)+�x�� �u�<���K�B��b��5`��2��lj.�L���%H� ߇t�h��ϻ����N��E��C��� gn}�xa �<$&��i���=O�D%&:���u�oen�'�ʠf�+�M�tm%�(���������ϸ�z�Z�o1�M&Y[E$ [���8D�#qML�c�O}���A�����ִ9�T�n�N��G�1���8�U�����f$��zǏ���_B��-ϘH��n��pY�s8��.��g �򤋈�v�J `��o[�T絊����n�6�,1��w`�
�� 㻒���ٱH;X����*�AM:�D{<�?�{~��S]��AdJ�&�J"�D�l���"f��n���2�u�dA f;��kez}�(��͹�e�놾y�>立�Yd�s4�_Q�a�aB'�����`[�r�FS���!h\��_�q����b���~jϨpc�����E�*V���Q�[�N٫��M��d��8��2��a޽���{�L���XO?��:-�R5[C�.��%g�=R�=X����	��"b�G��O��M;� ٫#�g���k�����C
)`n�NᆞS?��Ą[9�,\�)x��z�G�Et�H��KǢ��c ��y;4	������2�w9o����x�V��#-d	᝛X_:���g;��m���{�YGG~V�m�@�+���R��2�g��0|�����V�r�6�Q!��^Y��	��:P����L�4J���PH��4�1Nd(u'�}���;�)e�\��i��.�*�AVYv��%�*���볉�U��ko$�X�D��G]�l(;�5�(khHX�:%��yE�Y��j��B���k>�MLF�mBB�>^�;���F����Ȥ
���
1���[p��w�/�д>�)?pT�'{-5�Lҏ������/)k5=�6$h�2���l.�Vb���Q��Q�e�|����	�E2��{�i���Cɿ|�r��Nʭ��穾�]J-R���6�3����
���2�Ȱ � -^'�a�<a!�F�;�B�M�o$�͘���Mj�Tn���_��mdoz
��Y���-S ���Χ/ؙ��%���ZT�7]"@�ք��tiW�g.���/��ͷ
:oh�F�����C��B*�ytB�������q_����6��O�@�W���O�U��E�%���:x���ǘ
Ή~j?�A�u�k���wD�U]����i�"�Д4���!�ٽ:���Y�N�GK�Aw�E�^���:��U�$��!�u���P�є����r6*�㯳cZ���]�ׅ������|���{��8��H,��Eg*$r����IR"��y"
�nN�e�����4���'�a�sUH�0�7ʻ�Y=�ѡ�xi�yڈ'��'��_0�db��t�v�sݘ?�88�&\|ٗ�Su.4�>���?�i�����O3:�@"�f��]ʸ�d���>���Z���à{��'`ns}F�6]b���O:���f#[+랸�_c���@��L���!|����;����i�n�U/ם,J�3g��My���/��ˊ(��@1#j��R��$�����Wu��*&��0Pr�RL�<�5 %7�*`�h�yr�=�� S�@:�@��TEmW����ٍN��ŚVE��[Ń�4�0^I�߳g�,�.�r)%��ma�ڊ���+ԎhΣg��y�z����B�h�%�)��x�o).�`Wr�*���{
%@���fy��r�h��٦V3$�<��CJ��LoBe��Ffȶ�u%�߼��y�El��'��� È*F�A۷���5�B�8v�R�������SU2?_��v<
�a�Z��K�A�}��sĒ��'�/e�{�Ų|O7����@�/+���C��\[����"W�>s�4������ZQz�1�}y��⛎�F\�;�mT�Q����u�h�6�
*1s�.�҄�/�݌V�k����H_|��r]������������J���^�V�(ѧ ����p�� E_�Λ-`ޚ,�j�h��<��W]�I��09��ep�h�Z&�ߏG���w�t.?ڝ�LQ�D�U`�}(DR<�՝w���qK�����࿶2XC4�j��)s��4�de}���zt S���P����}���\�"�8�ƃTIQ�E�1���:*�������0�ZU�sH��*�rnZƣ�v;ޮ��Q9�d'?�2�[��Ьd�z��X����_�\K�eb��QcY2;0[���_�>�o��k�u���5��nZ%��������.9Q>ker�2�(&�2�t�,���\��G�UzrV>��h���B��Ţ:�;�G�Ѥ�3��=4	+��(���֦=H����]��Q{y��� p�> �A��`s�%�6���%y(��wѰ�Ay�<�ǧ���o~!mG�='�S�K���:v��jEp�<
,��Z�Fk�`[z���H>�<h���LM^����2
���=N�ϝ)�P�>f:��f�>�b�X�����<F���B`-�E17�bR�d'����=��5r���� "usY���=��ef�}��&z��Q�%;*6'��[��������:��MyH��LN:A�}8���Qʳ�y &qk��<ڐ5}��;�.��c&�Rv1�K�l 4I<,�.1 %�ߌ�# ��g2�*lrh�Z`̥��A��*S�����a��$�5���Z*�
��������yM��!F!�e��m����"��4/`N��Jy��E15�v��zs���3u��8^ҽch���EIR��d�:�l��±�������Zs�z�=�C&J�{����m��wb�}6��e
	�x �%]u�BO��]0��3�L�� +_��z�-=K��u��d�JW EƯq�GF�KSܽ��6Qn�o>��@,U�`	���f����H�g=�/�L]�]	{���p؉\^�nOc�y~]�iғ\�b���A@���y�Uen��v�<oo��ԔTI����O�-������d�E�]%��J����*
 u&G���~��ʥ�SQf�Qg�����K���ak����z2GԠ�$θ��$	Z�|�F5��p�/�U#Y����}ɬ���"a�^�J�`&�-Gź(�����vV�ʣ�L�����;Q0K<������Ŧ��L����)ԉBK��c��yVPZ"$�R��L������qojT��H�F�r�Ջ���{��G�iͰC\8}Gȡ�B]�s�fy���d�׮ I/�/Ւ� ~�v� ������yw���"pch8���w��ro�'P8���JRjaN�?�Ш4�ğ�z.]�t�<�Ҹ�`�1������W9��rh���/�aӼ�'"+Yke�$��<�qu��Z�Y�6qL��|C�����:4�A�s���7;ע�\��u]g�ȿr�[��8�aPz�e���Y��y"peR�V�s�Q�O8Q@ ��R{�,�����j/�!���PK1Λ�xE��+�d!�3i���[yF����]��8\����?�svmus빲�c2���I3�M�/������?�h�#���93��l���J�SXWs`a"����s]�����Sڿ�#7���8�ń�#p�)�#R�࿧����B�����PN���d&]�n��a�6	�p�u���eGU��}[2���R,���6Km;���D���Q%\��$��5�X7a�=�j+�}�+���Kz�A���z�i}�)�"�8n��+ڎQ��=��d�-䮼�h�*��d�UE��^%+��U���]�W��h$��ILآs@ƊDlyh���^�\�(����+�qJ�bF���w�D#-�܇��Q�n-1{1��CA�:��6d��`�\%�;��w,zG!l�8���
�W�"�ā;�F}�ˇ	�i��A.�I/�f����W�Υ�а]8��0]�H�|r��'hz�t������c�u�͒:� �!�)⟨5���L��t5�\1s��0�,�Sj~�۲��Qb�x��������=ނ��ְ�a����v/�u?���H�V�U1����Knn��tU��v�p~��\1�p����ж��c�զ��ߗ�WM�W�L��a��=�ܗL�
�At�A�q��v[��Za��vdhp���W��p����-���׎��F��$P���������E��(��{�e[��ۂ	�)�|� Vm�?C�xu�?��o�716�� z<.��B���GF����%v_����S��K���	bM�j�T27��K&����b2'R�כDf4�ݴ@���z>���1�����tl�/|Kx�A�`���	�
�$��Pf��	�3S�U�m��Vu��a&I�v	Y�6���>�2B�Y� e�@��J��~4Wy��/��6µ'i�F����`o���n�MS�+��S,P�^.9��Da��}l��羇Ef
�;���F_󇠫! ���^V�zS��}EX�[Q9�"��w��ā���)��cn���<���{�}tM'R��/���b��x5�lY^b�S�(���mUV������10�ʆ.��S����	������1�HŞ��	��L�ғ�F=Je���<:�m�	�`h��Z���5�m���k���q��E!��@������hm�MS�(p4��_��X�����נ��[�y������/�mm�T$ϋ��t�z?�A�ʜjӔ_Ԋ�d`��0']�q]�� ���~�XG]�b�\IɊ�{]e�#�đ��rS󮊨fjh �M=i<Q��8�A����Nז�s@�Y�3&�w`��wN��Y5|�y���x���Ђ���c�cz�5�(�5.ϊd���}��:Z�!-�o-8��H���i�^[��$�,5����@�Q�#�d����ɮ��@����L�x_<����j�(����c-�����(�w�YJ*��$FʠD��f��u��m']k`bed��R~��X�m���t�Dva;��:DK}��XS�F��<�9O��R-�F6��F>C6��'ԭ�d=3��-�	����;Jԧl�����sѪ����K�p�/.H%;���:qq��@y��-{�c��)I�'���úf����T���'y�?Gvl[�t�w����8�E-���)H������%�V�A&6���W���Z2"<���2����:�[���Zp2zϝ�{���.J��_�����d��81���?Wl��`W����iQ��ǂ�aB�~��;��ׁ(�T�W��y5�x�$G6e~����7�>w���; }�	��Sj��V��<>�0�u|5Ȍ|`�,"G�L9맶�ՉMB^L�Fx�kz�����x�W^J_���}1�w�)��l�1磘��pR����޳�&��H��`�-F
qݕ�P�b�E`�rd�a����z���5�|�������aŒrɞ([%/��3��&F{���о��5-)E�_@=���l���K��Ji��'�!�[g��??z���"S�hK���U�� �>�� ,Ȥ�O�;������xQ���,�YM�<�3Lb\~�F�j�2�S,�%���c�G��H�6$o��+Ҋx��:�=,}i�+�.���=�ƫ,�B��֘�V`A�D���4̴������?�5��Y��M�������S�:fT;�Z�z�ib�U� �-3��ub�L%S�������⹥յ0����"C�s'�*��<��w ����V@2Y}}�6�g)���6���x�oH���y�g���Fqh�pФ�U�Dc�O�S�C@�� |�t*\
c���Gf'�0�Eb�-%1~>O�^§m�l��+�\gX$�f���KR$R�S�aF�r�=߸�p %��*�>�w N��)N1�0�#�^Ks������D����zo=GѻR��4�2�gt?����k���\���P�#9���j��%�eΤ�Lln�Ү��^8���=���̃�5�%���(�2��a�n٬��!��k�4{Fs5��VQ�k�l�iiG�k�4E�:�����Ub��?�G�n93�����3%Tyt��b��o�N��z���7N��r����/�	�#��B��t���� LC�G}�3l�,��+X�y<�h�uhu��P�9�!L�����Ě�mt��P����ͩ�������5pe�o������d�փ�(����j�#4�W�˒/P�]�������a#�CH��hv�8��|���փ�8
א��0�+Pˠ�؝��W[�%��m[�d�@��4O��f���m���RxMZ���sR�4c	��V�Nd
������cu��(!��i~�����k*?xY�dM1�OjB��S$8,�u�ɩ�Ye�$	-,��'"�ڈdEu�qDԄeK��ӿ�Ԉ��>d�u2hw�1��A�m�j�S� ̧9� ��A�|M�t[!�<��B����Rx`V�U�%�!/�M�v�����x����Cȵn�`�Gl2�~����|�~*j�.�	��I����i"�Y���Z����c�2y�>�8nh�Q��{��l6x�`��N�8�q�Wõ|�f�/K�	�E�N�ܱY����BZ��C_B�����b��tR��
��eЁP����z��\��`W���r�čꓪi�t��/�	m@[#/\�Z�
��*�G�E��'h����v4^B-��"D�&v'=����]���Wq@\g7�,���b��VxF*e�I=��M"���f=�~);�S?�  ���
D��V����൛x��xTV����@͗P�{5&-�G?�_v `��������/�`��x�N{�o3��N���y�R�ⴰ$,��`x��Xq��9��3J���$�#��ZQ浾��(H^�o\� '&��ȃ��Qh'�I��l��E���f�Y3)ݮ殧�Ӽ?z����ҳ�@<�:Ag�.�� *�8��<F���{��옗��a��ڢ�����Lh ���Ն��Z,�g�!�k��j"�y%#�f����S�7Q�lTkO"չ�+�]D���ŹZ%���>��G��}\�a����y|Z�J  �1;��aB�1���
�]u�����M	�(�ܤ�"����l-s��Z�L�y:�e�>�zJe�6)W!�/��KjB3ǎf�V|�����s&���[?z�w5�[�%�+i����M��p��L�_���Cx��� r(�D|�F6͠j�cC:�Do�I&�S�?KP�19��Nv��H˗bٷή� �$��Oe�k�q9'A�j�>l����8g�y�R{ .��R=�8�+�|�3�.5��M;�(��ǯަ�M�0��/_WA(�U,�2��f�i^���3EF|��F�a�ֺ��z��S`kC �j�7��;n�]�3��bɃ��J���$d�ێ_SQ�bmsM�P&��b����}�!!��<�)��V݅��n��{��4�#*@%V�{]~�?�5�<#o?�ن����YIP��=�B�N��bn���}ѡ���\q�V���CZ�䇰ɕ�FL�"���md�A'�g*Ϛ����K�	������4z��Qq;w$�����|	�����[�K]�Wl\ ���$������60�U��>~+-�6��L'p�\�y�9f��'�!�B�(�)�]T���}܊�u�e���=�g��"b���jc�v��s��b="��a��ٯ���� �l
 /��_����.�}X�06u��? �d
b�PS9�4dL�^>��=�_E��XA�ՔE|�;=N���m7�/Pm�
>h ;�b�賵۴z�L��v6���_�^�(˨�
�PXjG/k�g.gʎ8 �C�,x��=�}�a� ���;��B�g �I٠��L(���g,�XV:r�7���ރ��l��,Z�AĻdt���MA�Q1�:{�w�%�} u��#��K���c$ma>]yz�E�_Q�	Hq�.��O �T��_�fDBfXGɛp��^ZYa5�gQz���K��{دxb �Y#��1��D���4����c��Ŀ�	��|ɶ�h�M��޴�O'e?���z�4b�%�~`����3�"f��������}:�3�L�̃�)���x|���C�rX\���Jg!N�M+�2b�O��R���-��x4S�i�chƑf�w8�.��f�[r0��e2�M�I�\]���y�-�a�O6�V1����"mږ��'Z����-�b|�;��]��m��*�4#��9֋��j(��p�]�� k��.J�����U-  �IP��@(W++�*z���+�c�"��N��-$&�O�����Ӯ�RGgIJ 6@���Hud�  �����U��o܀�FN���ݓ8����h�(\9|G[��w������s�T|Ŏ�Қ���Mh��e��x;�A:M��O��ߧ�/ �n��I��V�yB-�0Y^n?n,x��3���/�:Q�2�E��+�=F������4�w��I�]iM�c�Z�6L�=��	ȎL�H�AKM=��C���V�8�����I�p=�~5�ʸ>4F�.��J!Ԩ�}r!n)��;�~pA�z(�z��:I���N>������O�q���l]�֯
�P����Q�ŀ�T�L5,�;�"�Omt.���#g��c�ڷ���K��ax����0��Gȹ�+3R�Uq"����iL�H0Zqơ��t�2�2I&l��D0	���.���=r�%n�}�1QKJ��Gvء��Z���bh\��Pf�V�n%$��:,����ކo����b�z��nI�j�a-�4 �F���*�c�h���h�|8�j厌+�խY���xǈ��}~Y���y4�B��i�F�t�>����(v�� �f6n�e�$N�ޖ��t4ڗO ]�ٺb�|�����X��j���^ށ~Z��~P�<ݠ�[QlP��d��U8�,'޻�B� &0����0b`��WsZ���7����m�L@�	(��
���E �㢭�i���U�S>����H��JNP A$Y���7c"��Cϩ|�m�AjOP�\�H2��A�.�De��UדyN�J\7�.Ej���hb�:��?���Yp��5#Iƥ�8�mB���оZ�"ɤ[o,�0d� Mm�o#U^҅��?Ħ��j��IR����6FG*;<C�������M*�S��M	���4����||�ID�M y�i��;��F�X��A\��@L�ѷ�]���G[j�>��n���å��V�����%��y�{�|ם�aX��4_�;F��\������t�nj��)�hӇ�"M�B:�x��S�p�^+��!庂c�/��"T�&�Xm�$��:������(I3��"%����{�'���N�ꂠG�\j?X��0�C���w'Hq]ӑ��:�t��Jv�6/⏉�G��;d���Uy&���U����4lE���&��^R�s�שO*,G�6����4�G,�m#���1 ��Xӽ+��pW���ju� Ъ% '���
kF$�fŤ�x���˟%���;�{����{��i���]L��v�ziI�|�Zua�����SѮV}U�q�~|V��p������٫��P)Ժ?;G�{���Ve��T�9W�U�$G�Bӻڥ�@�m1�_�xK0EZ��k�,f���e�*�
'�~(-B'*5�񭦼Biv�E�'u���jل���Ú�w��k�9>��������i������i��)�Ι~n�t�x�N��M
��:��iXw-��Pv�m��'���w˩ЛK��l��J�7��:����b�؝��?QQ,K6^���]�_���g��-�����o���6��o�]r�'&�ʖ�YL쥏��lM����r�b�R��3�^D=�;��z
�쫹6���&6qyϴ��q��v8��f�+�� 3��'C��'�P�x8�Wٟ�sOEo���.n~MV�4 ����v,z����=�s�ݰvZ� ��B@�;n�#ci�����;��Ӡ����&
��!��E�Q���<�P�����.%Ћ��4�~� �,֒eM�=�׸{�Umk_�T�t4xK2�=��`
��=�k�Ԁ�I�Ai��ղ����ڈb��?�R�l�n������T�D�5��Jc�HxDQ,�
Ǣ���J�}�n��T8�h0���0�|�xc���mu�� �� T���g��~}�xCAe��A�w���L3����J����'9��-��@��F���1�[>G��΍:a.V�p��Z �<��sB����L٢a)B�9q��3��>�<BQ�+(����6kb��;��lq���rh��QS��0�ɮ[N`�y������K1!,nr(aG����^;�/(ZM�Yٺ�3�ה���w�s�w������b*YDf�}�;7^���~�):��d�3Q_���վ���D���oI؍��.��:�㬍�+�0�2�L���������Z�ETω��l�{�d��M0R>xXk�z>�
�-�Fh��E贼��e�����<�y���9��6�fL��~^=E� ��+e̠V�j�F/��]/(��cB�����i6:_%R�8^@#��͗;�䗊خ��1L�# �u�b����\���#���k"�+ͽ�jXy�b,k/�^�������BP�O�.0��'�e��!}SJ�bi>�*-3�����3*Ğ�=��eE�& ���gf���nދW��; Ϲk0:[ؓ£��Gq��2����yN���al[򟐽w'G/�Ť`���)�0T������"���:��39^^���r�7\�cm\��C�m�tW	���m,�Z������]��JQ?���C���
�c@�mb�d�e��!L�����-��o\=w��~VHB����b�u]w2�wlm��⛎�����es�t�߃U-�6�G���G�(�$O-�,Su�6g�v��t46n�en��{8i��郠�H"����^�f�� /Wa��4_�G?�M~eU�l�ڜ���vjه�`��͉h��:5��`��nL��NJ���/Qlq6сZ��O�Oh�*z&%�==��Ż����e�����K��t�'myW��Jf�
6G(��K.߷~�p#N��i|�T����V{��t��0�M3/�����^����n e"^����D�i�qt�f�����L��к��5�%�*�M$(l�l�=��[	����5F��Ix��_�bh�`-�3M��K�A'�u��%s��&���ku����g7K���_�-X
�K�_����?ή�&���[��	�c3#N����WK���[�׽�F�<��z�\a��Kj����v��3�|�Z{���7Ǎ�o,�'���N�M2�y�a,�bD펗�� Mڸ�v�G5�ۂ��C���eW'A|�ݩ0isԏ<%W��?o�w�Ӗ�E3yɓ���WR���qw#�m��$�'~�&iR����|���G��R�
�R6'G��{O+_R��H��*��#��{�s�%��?�p���;��ַC���Ӽ�vN��V����rE���b����jsD[x�U�_h�w�*f����̭�F�������&����mb^�-����t�;
�A�M*���`3(��w
�!�Nێvx`�c��'��G[��ψ���O�^g���w�, ��Ǚ�1���v��zhK2����5j�����8 �ڧ";<_������8�UJ��,��h��ڱd�vQ�"�z����|,R�w�pt�{�y!~����]��28b9�	ܙ
^.����������юx8O��'�{�xJ�d����gC�?}c�\'p�{�d}�|3w6��jr�`����xak�/U�qh�Bpڪ��Ƥ���'��wV1���+R��^S�G�$��RM��2tD�e��`:���{f7��'��z#izp��yn����!7@'O]Z��9 v�h�`�R�f��8")�P�vM�*؊l�jfg21^O��.n�]��@T� �J��őKk^����V�+�_#0g��5#P
錇�cl��k!5s`"��|I@KC���Qʖy�]�����q�,��D+�xE�%`p	j��f'�
����
���~K3�\�Bm/�;
YӲ��04~(��KE`!ʮ96��92I o�d�շ��}�WW�|k)�Z��x5y�_�-=��=������n7�YT*���=�!f'x�}�=힔�Pg�4�@���"���
z�=:�Z4t�R�Ο.Eu�#/F~�SL�94��N�C�H\��zlPR0 /��G)ײv4�A�GMk����E��*�����I�u�&���B�� N�?��ލc��-�m�^��e��~<���"�SQ��y=�9�BoÞN��r<_����6x��_���lp��rU�N������n ?�G*�gE�����P��=N��/ҲDс {F9lmH��I<�0�z���"����c��(z\�`]`$(��g@��A��#��k�$�Z���)�A���=�8�f���Yb���$E��/4qB2ב�pOQL�&�|&�'�{����UG�J�!�۸'|�5Ѧ�‴��Qb�PE����-]C���Q!���?��y�@	Ell4{2ɽ�ʮP��c�H�����u'l5.Rթ!�'��9>�s?�����r%wΡ�%��%L�z �Ǎx�\�6�QTѓh�h��7eS������O��G��$9c�q���B���t� �3�n�Q\����́���%�׀�77UO��{˻�/h�'�P��o*{���PpA�f6Wyњ�(�Dװzq`:������ �a�,��k��<|,���--�5�2 H�O[��/���ѹd�/�G"N!��G�^y-��e�)�����W�Z�Y�m\�y�95���w�R&: �4��FV�x���d˞�4ƶ��`�,h��E��ҿ�ɯi���i��gQ++C�\
x��6}?4)��I��-�zuH2B�P�!%A=�b�>�n�ly�hK�����R��HO7���C®w1e����¼j�VH_���C/,�i�sJ�T\���{_�.��[�e������mCz	Y�u �wH�&S��x�z�x��Om��7` �O�f���']�)G�i�}���/��>�E��%X����"�N�8S�Y�x����(w��bO����0HR���|�H7�څ�M7�=�[x�$����H�I
m��#��D=1��'3S.��'dq�N�l���8���Fʆ��uG���@��+�,I�v����ft##l>}պ���0BU��9��j����
uQ ���:k��v�����왤濼^��)G#=�؝so�I'���PW�^V��뀵K�Oj��_͈�?����_�
Ȩ ��T�K�k~woOles�Π̒G�\ G��^LS��oӘ�d>��~������T[?�w�q* ���M_����}ہ�y_ɢ�A�_�*ePV�)ݯ�ܬ�oЌ!��LB��״2*�,^ �a+���}�ɩh%���xG*�=�3��.? Pn���0�5�VWP�m]���E���T��H_��Q�)�h�ܗ%�xsK>����d#�N�z�֌j���<rNl�AY�2е�&:?�j4.�-o�3��n��uW'Y�~�'y���B۶�!q|�V�ϧ�9�k5�쨈��*C�U �&l�|Z��/��1sc�Vʈq^�|��e�':��t�T�Ι7x����j�^aueq�]0-\���`�d7���ˇ̈�<�[L��`2p��a���T�q���wvC�0�gtw ���ȭ��	�Y9L`D���I���A�q;>��7�u��7"�g���;��Q��h����-잯���ܟt����-��o�'A�i�(����1�e�u����:�uٳ���m���\�/��p����l�N	��=��N#��W;hxڳ�EA�k�R�`����Q�s㇇kf<����P[y�B�EL!�+�}�T��ع�6.C�q҃o��S��d�RoS 	�)�˒�3PŠ�a��D�'�,q`�mʌ��1�T�E3�'��ܛ�Ak� ���jWe�Zw�T<���z6�����0��޶����n;�����sD�}o�,K����Ƚ\6;x�6^�6I7*X�{�zDP4x��8>���ǂ%�N?�vz��Dﱂ��Nk��I�݌��:k�g����ͷ�ߋ��n���b����dD0�~`��i��s��F�%߿��3�S�
����SC�2���E�4�d;���̥>�����F��
=c�㎞#����q.��$=�Ԇ�Ψ�=NBe��#N?�?���[�m/��U�cc��-v=U��;�}!��1�=xJ������\fx��[k�2�aݿXOfN��(S��4�J����14��!���A���e���Y�61���4_�ӓ�|ynUݹ���l��(��k�W�"Fv�"˳ (�O���ίnZ?��/a��t,�v+��S��ɳ����D0����u�=j�E9�y*�uU�����9���#����^ԗ)�"�`-X�|_����W�br2�N�[��Z|'wwL�)����D�����e����Է�<�����u�*���`���ƣP�GU����&<`�r8�Y?F3-|���&ڲۛ�s�䚺���1���;o�n`���iӥ���X�b�؞Mo��~�Y�Iу�w��p�q���b���r�=>�8�H�>��s���z�.�>8E�2]{I�d_3=��/혽8��	`����Yh��4=tѪ�/]���g�P����6U�lQ����r�L�0��H<�@���!+�&Em��)� ������j� �JUП��Jt陫2��e��B�{��x��
�|0w�V~��YD����I��G�,"���Ke{�3���p*lJ94�?�ט��9	ڪL�tp��"<q��I� U��������qo�-�MY���[]r��TNPG�
5���ޜk�A9���~��u�b0!��]݅Q%����8��#;�-��gH	hb�j�Ke�����������Y���,�Lw�1�C6*KW��}�l���22J ��s�� o��WF����k����q^Lr�iy�)���I�l�� ���f���5�1�!��m�-<CAJ��<�m�/�0e� ���cȵ�Qt|�j��	]���K(�C-�����{�@AP�*�����)�{�V`n�a������g92}�_s��P��E��E�v `7�̦�p�bz��1?O=�:�4�n������W�iq$��H�%c�3sܨ�qC~~��xB��K��v ��ʇ�BVƐ��*��d�1���ar�0���_W��'TH�N-���z���U�5���Z��Hc�S�  �[z��B��%@�Jh���ڪ��#v>X2�p>|Qq�V V�T�,Rx���"n���$iV�Qq�}e��tѡp�����7"�����R���^1s��V��n�Uv����O�r�;RvAL�v]�K��e�4�O�ZЊkQ��<�0j�����l�g_�BhB;�A}�Y���|05��ZZ�ݮ>.��8��P&��]f.����aNbT^s����yR��l��D_��!Z��5g�G����cM�{����F��s�A�ōr��_iK�~��~O�3#��7�'W�,�}Oq���u|oʙ�@E���y!Y)^�<�]�� ���DKE���-�@�]K}�=1�ίf*{��5����qL�=<�鲴��G��{�p(����e5%���/�
����a
�=n@���Ċy:����'��EK�I7b�k��G�����j���ɦ��:G��_?+�B�J*b�m���q�۠��ͳH�U��	t4�p��F{��B��|�B_FVէV�:�YX���h����'y�K蓈�O�⬰��1& �Cy�^���hB>g�5�gN�8�V��ޠ�_�ڧl�n�_	�d��A.u�b��lw���̀�����J*����W����Cjmܭ���?lژ�FC�i�щ�A}�% �8C`+��J>�tu��E��U��%���S��Y���3��5i�W�<���t�2,�2Y3B�Dz�/s����ܯ�P����DH�t��2�.��s5����C���I��[c����Z�r��"���Nd�!��+;7�������uR��xf���{Y��ڡ�����!)3 ƀ��B>��&y��Z������
��6��[J�nʬ�p�*��#�i��N����j=��5aAE�!�����z�2�����:
,c��2҂��AL��J��k��pCa�D�Q�][��e�$,"��;�q��U1`���V�z\!�ٶ9~\\_��uxƅ��u��Ie�@����u��3��ӷ�۬�PI؂�邀R�Ar����I��k��Ir�����vV��e�&�+�\Χ��\�,o�qVǄ��&�k�q�������޷_p�`�_�G��p��Iۯ"��_5���������U"���pX�� [?Ia���O9�	���)��]Iu�^��2C���G��dj� ��p�����3\�eJT���aXw�sb׍\.=���(�c�w�P����3�|��;ʽ*T�}jd��2o�i�5��`����^krw��yZ��~�j�Y;g{�'�V�����߃�#���o��%�	0vǧ~cg�Ah^�UdQ�G��J�s*zo��R�sCĢ\6%�M�񿐦��,�F�wWs�Q���~�V.ӣ���w:�{���ԡ:���m�n�\�O��|~{�j/Hg}��1�+��'b��1%U���%���.���c`�S_㎩J���;M̄v�} �+���2P�M�>�ӗ�	\i9xl�ے�������\�n�S�m��]��<�IM���glېA�2F�јО��(3+֡�p\��H&Ʃ���x�dw? V�`a��@ڢ�k!�-+$�E&��U;��4?�ß��h��=��l���\<�,k7�_�Uy���"�?�I�������ǳ �1�j0�\K���Օ��(T��A��̈�IMZF����;7#�f�I�6�F��m��e{L"�l�6I��fl'me���$��+i�r�]3���IB�˭<��|�-� ��'G�)�ü��C���Su�J����k��|�d�x�g�&J�Ms:�x��ڴjR/��&�ֵ�{���]�ܒ ���h����˅��8,R`U��
(Vx��Ho��r��}M�7�</�M�q�8�[���ճ��,9�02�j��*�Y��jx\��_��̾�����j޲#���#vD���Ō�jwI�n2���C.�ec6�����T��p�*��Hd��x8dZ�k��$ͩ��g��#�}���WRԔ��4@�����
#���2<��v�b�@��U��������������h��(Ԛ�4�_bG��ь���,�ƣ�ګ��Kh�7�4��Hh�_w�d.�q�N��9Æ����hdt�v2GƷw�������n8CI�!��O�P
\�J`ܨ{�O/\mf�(��u����j-�x "I�U�Dq��tῴ�7�UF���4�l��y�6��n�����	�V�Xƍ��<�WM�v��$O��N��(����Λc+��}/x�&l��i|��g/ȣ$��!�'��yӖ���|nל�bX)P�/f��2��J���|,��2�Q����#z޺d��y�&y7C�a4�;>b��=[��򿜣���o��җU� �[W��;����pjэf�X]�C:�}���s��j@�RΤ���:��7�l�l���ܹ��V�Z7$�Nx�K�N1�cu(_������q�I|�)<���r����{9�����Tss���K�i`��&��ov>�2��#iY8��WI������'zhهW��L=/�*��]n�Pd�V��e�}�i]�V�y���-���3�B�������	3IU����r�E�T^�bk���s9�蠈��v~�=w\�KG+�&m�X��P�=
*=g��o��	��vC��ы��rL�Dz�Q���6���.�?GL��o�\��?p��p����"���gP��1�:��/o p|��rr�6�nq�h���bx�y"�6���ȸ����܇�[Қ$v�C�-�$���㞐�PW oA=�k���u��p�n1O�ݝ.�i�Bk��rG�?��9�
�ej��{b�@$��>�����񃸔����s�~HĒo@@Fd�H�5Y��X �����)W3X@cr尤��;2��jEK����� ����;8� ^/D=X�o�C6���}m�q����4/L�}Hw�@�}�����W����+���$OՄ��4Fp�c`d�<�t�}�BF���"mO�9H���kQ�jH�����d�ϼ���G?C��p�M�v�
#�z��op�`��J%��P�����K�a3�~�*���hq8m���1$���>)��b��C����(;��U�;z�����,��x�:(û��.�����8��׏X@Ǟ����W[>?����m����y�p��>��$�Q�[G��`��B��uS�<j����ƫ�~�Qۄ����w
�*lY6�:��P�{�(%mI6�M���_�gv3�7z(<�wb����iI���<�����XD�g��ݣ� �F�%&� ��#'�)8�W� �c�"���γ.`�ŵ}s�{�v[�'�!�^���o8I\dpke���2���<��H���6��iP��-%�;n�GGc ���j�ȉ�dצ�옴ۢT��	�"H5�JЄ���VW ���8O�F:��f����sZ�@��HxV�{A��Rr+H�E"s�� �BY!�m= {�׿U6�!p�j>��e�|P�.Ǭ�+�\x�,lP�>��@����rSl�x_g�co��;&���?��-����i
���ޠ>�K�N'
�A��S�	ib��9r�s4c�8�4U���A����gn���ٲ\_��=�UE}��U�ڕ��,�Ѣ�N`-��k�[;����F�F��Pb��QUC��a�05S2G���Y��s�$�����F���o�R	��=��4�,{dG{[�3v�1�"�T�T�Y��z����'@���J��Z��z�ǧ4J���މJX�����������������+P�'���O��`6������Xi'�L�(��<�v��b������gP�S�9���x����ց��i��0xH�>ۦF��AE�ٵ�Cn��IqHw$��Z���U<�����oH��ڵ�.ޗ�h��=�$��GTeָ,�3�a#bL�^͘\Bpq��<[��z����o��.Ԑ���U�{
�Wīp֬�*�6����p��/��t��Vϴ}k���܇6���;�H�� ۋݑl<�D�q�5���/:��S�66�: �r�I����6H���Jz���\Ր{<j$H��T��f���o����%ב��A~��l���j�(Q�Fbn�`�T��V�Y~��	��Ͳ�e"�Qs؈�Fa��M�CT:���J�P.y��f�1�x��� M"��͛�Ɋc��mE�:�K��4t{W�-b�"�����àdn%k���d��a�;?����ք_�&:�A�rP��ir������P� �e���f5ҿ
�d]y$��#5��pyE���A\߫h(��=G{	F��aw�c��*�-ő#�X��?�T��+|b#?g?�̍���Iȗ�ܡ�
�s2΁tP�>�ji���L ��K����: ��֣�^F����Y�1E4��K(�Fu����m���7��.(\87�%��-
��k)J���-o[��3��i�.�{�?���20ky�w�Ơ1�%��N�c9o,(u�%��7���*�"ے}���$�0��>�,��`i]�k��F�?J�=����gU����0
UB�����e3�r��G����Wt�W��B��g�<k�u�j��gxwo^�@?|i�4d!r)��j9o��3�&[�o�ov��i-���&7��;�܊�[���;�����Ǖ�'���Hf��7 y�Q�ʕ��X^2�&K������C[X��y�B�.�v0�����De
 �N�mw�sn�?2�
���"c��^He��	H��w����h!���].jP�k��,����F�8����S=�ǮbA<��S��iK_�6���T3�Y}�L���4�}�lq6v�.m=� �B�ӪG�>a2��iړ�����$HaB��]PH��φ��7䯧��Õ���8Xl��x�j��"z�lp6�y��g?D|4�.y��h�U�e����A)E*�m��#*O�?�cF	����̓�n�
�Q�p�'�~iUL����a�����x%��BV�I�D��e�Ր4{
�!�m��g*"�i���PćΘX�eȐ�h��=�r�$��c뉿�)��B��>��2�S�Tc_���ذs�F-Y�!r���pNE���,Xޮ[#jU��QGN�Pt (��W��Ÿ���ɩ�;~��T}R@拺ut�W^'vr���D�X��f�2�zi�[��q�4���\��6����M�p����L��C�x,���QLB(�������@�$��Rݪ Vۻ����%��͕��(�#<ox�E0	V�ȣ��'���ɖ|4���j�g�b����󤩑q�*ҔYeT�r$	��7R'����dT�����'!���%��s�g4��r@R�,˽��F����i��r
(�\{����gq�F�;��G����G�|
-z��5NN��AT�p8ꅰQEm�'������o�/U�0'�%Z�����%V���/�{.�� ��o����� ��$�r@�r��8>��7�Wt�����!�TǄ9>Ut��bx��9Bd=�e�2t�g�`�1M!
�Q�pX,�1�}ߺڔ�qOӇ^?������٦>���0/R�ai�� ��b���1�m�%Fu�Y��/�5Ke�]�I��s�I5�(ʨD���m�?e��"8�+Pk�c�S1ib�y��+���%Г��d�w���㶔����]�%�}�j��2��E������]Dc ������$�>�ҕm�d��R<ͽ�xuo����yj��v�2��RCf ��U�}B��fr���[߯ŉ��EJ����Dz�Lc�k=�p�����Sѝ��
.+φ{
�|��8�e.���
1�~�J�5nޖ.y-��E��N�Ab������᧍��q��P�h�P�w,����Ad���^KFw5Y̠��G��k�T3+�%�X2�����隱�� ��6�.�"˜�� ���F���W��A��M��ߌ�bp��� �)��_P��edD�/sᗠ#*���턐�6.����Oնq��G�ػPw��J ���(��R�P���(M�n�ʢƤ��/���~��*J�u��Y!:��vl.i�ᚍ`kSB1*D�5�q)����p7*��*S] �3'�lfNF�bcZO�%j��(C���ê��N$d�I��4��ǘ���6K���M�{���׶��T�R�יj��U8=�W�M�Wt�/�`�m�!̦t@m�5�7�~���7��֘�O1D�%����o�*�L�������e�Z����������bi�/�P��ꑼO�X3j��ghV�ؓ�hdo�l��@���֓
�R�V��ҵ����3-D2�T���􏘺��TA֑�r̒.������=�dF*�S�RYU6�V{��&�b��<8�h�-�	��m�F-�>;�u�!������3���r)<y�pV�N��n�3�8����z��'�)��9W�:;H�+�������f�[�g�+'U_V���ĺ�d��Y�e>�BIԙ�*���������"��}�L�$u�d�(���������<X;H�A��J�6M1� J֗Q�Y��O��H�:��V�w[I��K&��x���)@�"�qVF�� &)���Z�r\z�-g8�}����o��^��q�x��^��v�	C�ZO�e�gwl��[�i�����V7o�R~e������M�hѷe�Y�N���6��DUt��y{��5����k2��e���~Wr����au�H�K3+�|=����y�n1o`q�ĬfxD����S�Cf�y$���8�>1U�L��u������-|[�!ݕh�9��I�%!�I8�m֣��1Mh���"@�����%�:�L�ۡ;���?~6��7U���aH_�$�^�a���?�,�.;}ٺ"�����U���	<4�t��A�_0H<UAF`h�mn +���*r05�<�R�,�mkر�*cG�X���[��������4�[�:��=
��9'FH�ش�acw��TN������"%�o������r�>�;�?�Ǉ� �V���I�����f��|�#�⭘��`>k�e�otQ��D��P����I'J��_��%�`~
M�`�6�(!���9���&Dze�h��s3��������FE�% �㨎�-_c�{��N��<����\;d���a]�ܺ4Ų @�\V#xq�B"�F����}���wDYF�$B@���t�x����#/�]�hsqТ~��bHo�K�]��/S�_բ��"O�='�+�����"�/�w���l*{���2��|��"0O�f��h�md	��v�?��q��[kޯ|]G�X���H�.zN�S^!��Y�kS�՛u �h^gyO�d!\�&�tخP��0�!x0�����\�0�H��M��1JDع��g�)�h�_���w�	1X�N��gi����Eٴ���߲z�A�D(��^�Bj�;��@A���쉝M���n\�p�H��ON{H��EQDa V��� *ZhWc�k�AK�K^��A�j��G���A5��`�?0'x�����.~ւ�[�/����\��8�C��89>N�����zr�7���L;8��)����Չ����>%扉;*g��;��k'¢��][� 8��3i0�%A����h�^Ŧ�D��Z¸�?^���4����6уx�*��a���vT�h����/��O��Ș 9~v<�X�;���uf#��Z�R��E=�c�q�R�ܴ?5Nhy󫫱��pg��đ�@]U�_��@�d"1U�Y+Q����d �sʙvIC��<C���� =���-R�{4�ƕ��h#�4�
�x��H)5#8jI��b~��<&�hoqC@����9��T
qNb��m��=$��F|���B��d��R�N"��*�$Iq�p޳��T��+��lcEr-��(����=�VS;4�ܜa�YHU�>P�eR�7�F<l���`�҂U2�a$"�����[J��,
ݞ�d�<�;�ۯp�!��q�@!J0s�׆�>N*eaR@q�������;��#�AlE��9��d{�/h/�j�ld\_ <�[y��{B�0[rq��ao-����uF��Ǖ��$:�w3;�����*=�.-wɊ�@�}�����>�a�wO/����F�ⷒ%,���*�)�)���%	��edBR���u�_&�$q�7/�U��2]�3DJ��g0��;��#v9��m9�\`gT~~8��e���.�#Ҹ��b���R�t[�ҭv�!S��'��O�YO��0��p�r�kcTT�D�Eʻ��1:n�ӣ%�XMX*3�Xa�3��:��N�����toAH�y�Xm�f���scl�L?!�T����Y�C���p�tb#�]�{Q�	9r�l3A��>�� �Ͱ���Ϛ��ﳘW���ٸS|+��7ͨ��3c��;�Ȏ�n���K�)����ˠ"C��"���З��?�7�I����B�*56��(��ij���A�MH)X���e�"��Bf��)��� h�wJ;��o�ga���x￿�Ȧ,Žy�f�5�O��̂���o�z)���G�S�A�X��Fήp��K1�һ�;c�Z�
��O?~�tK���D}_^����%uו��'��Yrt�΍���:��R2A�0u��yB�>�Wv� ƌLw��� ��o�>�D������nM�лP�7~@�抡r��B�.P{�컉c��>�;��9�W�v� ��y�-��l%�"��l �K�`�(C��0��ݲi��L�|��Ut�e�$�I�ۍxb�b"� �������̗���t:m��Giv���r�-������g��qC�����u�i9�~�Λ��@�E�w��kc�mзr'H[$�D�c��CA���/�'�{ɏ���+�fF&����9�.�d�)�j���L�o(����hUJR��AZ%��ӱ���2��K��v�����|����c��m/��Z�TG�ܨ��sU��I{-Iy��B.^�ޯH�KRfM��Lk�=�3�'����e�w��V����xn̒5�C��������_����9 }�_�&������&�j_&[���3�U_�v��9��K������a��ᐁ�N�#G�E=�]��@�Kud��Тh[�(��
l�˵8>�{��}�h���R����χ۽N��3�ah$��/�D]�J�s:&%���V���@.H�W���i���&Nu�L�h�#n��+k�9�(�@�
�E�2��'Q��w:$��AL_A�.,���&�U%"�좐�j�����K�Mx]D	<��l�aZ�<������_�i~�T�_��a����nz ����,�;�t�zDQ�j^�U�E."h��pTrDӎ/i���Jo�� ��S���zCXZ���R$�!�_�q��(��x1!�����La°���/ȈB^Jݜ�T`�|V�X�j�:�4o���f���˘T�{�+��m�~;�U�n�ߟ��- ah�'�M��ac�����T��@I����2��"MSV�*�h�C��@�|��A�);��y������ΰ��剠dꄎ�v��ן\��`x�7u��t�;Tui򵒬3������n�>�� ���>���O)�?�	�|�O�$���Q)_ì��j�`�syK���u W���=6�����^�
*��/��	їp�n֊�����0+M893�`�/|���TZ2�y^@uuL`}hR���5�-ʌ}�9��HsH��a���$3�*��9������`�r*�<�o�6�ơ�/V\-�7��W�����0�+�H�پ���5̽@�	,��/����OѸ�gM�$�176�"�w���r���J�T�e��rx�(D���g�n�� ��`���OdQ
�{�]�!v1�Lto5.�Z�':�VR2�^E�j�^Q/H��vM�}�x��hk�Y�Kh�M�<� �|h��A%x!��Z�ꯆO�o����q�9�Y܈$�f��X��� ���OyzEx����u�;�t�:�[�!�������'0��Յ"���u1	:�J謲mv����^+��g�;r���C_�|��
�|*,���_�=f-U^r'�zb�vV��n���te?�	���yEo �� �d�>�P�5�{s0~P�Ny#";���:�)=�H�o\s��M�;+��.����}H�?��}eiZR��O_��	�j��ts6"����lB�l-Μ���?��Oۇ�^�\�e������S+y���[���]�|��T�����`}���L\�c��#=X��ܶ/ӯzڹep��U�T���D#�`U3�Z�[ڈ@���_�0�S<� 	!򩁤"N!��+%�`�{[r�� 1��gDx�He//t-ʹ}q>�؂�=�Ƙ5Pe�/��4|3.�������V1*���F����}��B�J�yY���j������GpBR�E�ۤ;yw��\d&f%�ٯPj;�w��43�oP��;E}�� ���;/b3tF� GI���o�����X�ܩ�w�A����5������JX��ͬ��xj��qx�#y� �,�¯����H?�(��R�6�m��MA$���ݐ0��=��v��(b��޽��>�}��QK��}�d���\L�"�2m�����ӰC�<o�\� ��h'.��|m�̢[h����p��U���k��vB{��Dq����H(`�,�7֗��溤�0�0y<p5:!G�6����)�s�G����R�3W"�9�o	��Z�,+]��;ޤ�FO Tb��@ߏ6�6�Zg�t���
I,�owܶI�$.��L�in,Zg/�L������5�2o|]N�r�Q�|4�����=�|���)�T����h�\�w���)�x���6܌&��Z3�]�o�Ahv�wh���hX�-c�j�����h�1�J#�Mip5���}�e�z����^�T���r�1����ə�i��~�zl�3�8��?8G����r���7�[���4;�TV��oG)���;�}?�g�J��Ve����l"������l4�b� ��6�,ٵ�r��Z%�g
S=bua����aA�\�5vk��s���9F�}_�4r��:4���𒤏]YY��n.�Qz��pG����) t�8�G�k�>a�#ܾl��Ċ�uyO�*�ٲ²�F�ڶ̤Ȑ���y5�V:��^��}���"?�W�-mR���CM�T���'���O��C�Se���4+�^�Xa�E��F��u���mʓ���ͪ�u�w� ն��^6pk�E��웏�qT�J*Z/��R�g{��ix���ò�'��[/YL�v�Y?(���A�&�J"�Bg�Y���C�<S�n��_�/�ai�CH+;�~dQ��-$	:��0�3y��s<�=����B>��op31*��@@k�^o��D|U������(J����Eo[�-���q�7��o��Q�9\�LC�U+��t�z���A	�>�Gj��E���l%��,w}��M	7G53�o��s-�_�/d���`��d�i�xf�w��t�Oq�������3��W��̷Qy�j�T�@�Y������
�+�/R��P,�#�]�g�\͍-'�~8Rؿ�z��:K�^̭磻�W���%�i��rte��C�x<"\��_�����n�ٕ��1ϐ�Hb�g���L�U�z�^�G���\�/K#A��,�F�<E'%i:���N��2y;�_�r��m�����0/޿1묄�Q��7mVO.�Ԑ��kG��`~�%�N���(V�u��ņI>[��.Ev�5T�WwR��/� P��,�h�C���9��+�m��pQ���
D��پs,M��o���x��`�}�b��M�?�7`��rMA!h���9	��j7,�{?1�@�����*M���&rǷ<͚���Q���mAa.�ݝ�v��Z_������g���O)t�(P稨������`EZy��w ���`�거ɕ>�"�X�9��х�x��=�Ԭ���+=�3 ��<��R�ν�2S������M��2a����h�3cÉ;�L�Rq���d1<����}��7�NO�!��t=6Br����?��6���/�N�!�O��T8%7��T�������[�f(��C%��bG �a���a��q�/��y��ۉ��ɠ��v�~���J2��j`�S4��J��]P�M�B��#q6�E�gI�1gK���K��m�9��"��83e�Qp�Iz�shV���5V�/�,qX~5��X���^�A�z��~q�+3�1����v v^���|n�Њ���~k�:�͗*Y�w���r�d�87dt�,3x��[�o��>�~[�Xߴ�W�/y�d#�l_-d�����^�6g.8�`|g��6PX�ϩ����P���+��̄f�yG��P������$�9�p�Z@A�xMe:;�"��ф��I���&R�F=[�p��@}K�E1�E1s �f��gRNq�G<d�"�}E�3]�4�:�=c���č=��6Dzg@��u�JJ�������UӖ�4�;5��/�S�<�`K\߿�=��Ax���l�H�L�Ī�	��3�D�оen���1�DC����.�Gc�d�����%\�Ȫ►������`���gt%��q3#�\�q�
W8Ô[��R�N�<Q�S���t�J��`,����� �*W�
[�Iqԋ<�"sq�߾"�h�b�zH��Xg4
5�A-@f���-k��q2�miV
�TN�P?^X���?�;a	��"	]f�G��}+R��U�C��dk6%I���8��g���8K89U�J���1i�Tp��v����\+~��'J~�Vnc�����ٵ�U��?5�+Q�^���Q��	t��d�q��I��jϨ����y�g����^�Aŗ���2�<c����Gl�C�	�P`�`���!���������5T/*<#�Vu���j͕ĄF��U$��\��t��I�T6e0���'w��^:�d�ɶA���]�0W����������2�0��Μ��m�\m�D��An�]�zм$x�
��WV�QA�p��$��Qv�X8z�xi��)	��T�M�?*��e�n<��m��m��Wzw��$�&�]�˦�+�V#���5/2�ɦ)(<j����zvkI��J-g��D�+���x���_�q�#j���p���D �R��\��oi��+R��zs���`���VrG��ߓ�,δ*��.HC��Ҩ��gj���i+�#e�����A�{r��z�:ȰV+��!����;�w����m�W߮�{`J���6j��X�I0.�n�ߵ��RBQ�U�#�:�	�ӊQ��M�"+����Y�>�j�o�XxB��%�fs�c"��\�C+f�Ҷ�i�wqx��1w�#S��Ď��*�+�D�E#��O`�����ѵ	9|LEn�Cq��s�����.Ѯ:vѿ^Ć�d��n������級	oզ�G��-�NXrR�f"A��K�l��cfa��u?CQ���$1�~�!��p�-q�(2����F��0�O�;ء���~��{&�
��
��6DV���E����u���� Oꌐ��ب���)��x�j��g&1h2�g8��hB���l��e^�m��@���Qt����,�|��sf�B	�u=ڏά�z�7��q�;s��Z{�Q�~i���	��^dQ-�\�*��Em��j�8�J�m�g�ڕ�L��`�G mY"E�~ޚ�BRFz0d��|�@�����iqj!|f�P�'�|��%�p��#��B�������R��A��n�/�d$�9k��76�m�o��L�!��n�*�oT'i`K9�p�1Uh�^#����;�w3.7�ϱ.J����n�(�L��{_?B�׀�?�R����[4Ƃ����g������n��E/D��rK�/�%ywï^.��]��"3�G<B�i�.��G�ccDᑱ��j�de<�����'zC��gx=�C�c� 4��#��ͩ�YW�3���A���BRNr��	�ܵ������M��LVi�������yjhR��ˉ��q�tܞI�L	ٗ(�����4+��Ղ�ɫ�,j!�ch�	���!��r��*Yi�.bNY�=��V��T�	a�'j�_��7nk�6Ȋ�Wg��ਿ�fL��-�)(;�w<�}*N���y"�n115'�p:����ky�t��I.dR�Ĕ��0��G�^V�}�/8=�N �)�]�'��ߝA8*�-�ח=��&u��y��Z#�*�5Hu3u�$}�k��&[
��*;�#E_�L5��X�����Q�ۭ�%,&�(W�	��7G'��$�#�	�3���(;s�z�Q���d�%���؜I/�?�d^t�YO�d�}�:�'{��L�K�7�=�YtyN�m�_�ȯ4������5cq�B;%U�")l!:�c0BYh��\S��IG�Ô���%5�X�as"/+�����2�N�{��+t��5�
���=��f
�JO�B�֬3�Ɏ!�N
��R���|%u�5x<r�q�u������!���!2�h�v���j`��R���N���GᇰM�*̐�����QZ�ܹ���dS|�lD�U��og辉�?f���sθ��' ά��l���i�Y�� ��
���ܭA����|q�h�S����p����
P��_� �V�n�0*�I�\�&���4�Q?�'v!�Ncc��f s}����R ��|8s00����vAI���k�Q�����2c�K��F���i��%=����F�� �uW��h�'T��WgUVp��v2$�*XP�.�1onx.|�7Ez�h��4=�~m#�z%��:۾��w���_V}�N���9O��
T��rec�#�Q- �#u�tU��ݑ#N@�d�[�W.H�@u�'n�T�#��&}��6}r�x�Z����a��r��k�g��s�T��[��D�s���8N�v��,����펕���>wjh���eK��q!��$͵#��� ,�ίb��5Kβ7W1����T�[kˇ���a��R�m�Ւ�k����~y��-I�}Ͱ����x}��2��d	�V7�;�2���� �X#��V�K��L��0�Q��?�{�4`�"�|���v������2J_8Fl�˵��e47C
�"���͞d!Q��7=n+^�Y���mD��$n����⒣���!:9y��b(f����ؙ4�̺Z�%QԷ�T~�JM��q;5t��R��y���]`�$xw3A(=�/���� �5�b�=���?@���z��T�P6�W�� ��8�V�,�\�]P i8�[�Կ�ڤ'8�������:A`#ׂ�ٹ0ƈ�[�F�^���8ΣJ|��t#�e	 '>m=�Թ4��5h��K�f�z����s�E?Kn��յ  ����L�ɠ� ى�(d�S�_(�zo��!I��r�IY͘/ك�/���]�@���C���гneZ��}dK7fuzpFC��7���/�K�M�ͽp�2X�k�-��~D�>�'�/�¿�Q��oL�ic7Zq{�_���_�-Tj[��B���'.�����JV�n���<���'����$C\�9�s����A�ZT6�l�]5�%Uo��Y�Ӯ:��@�Ĉ���U�X��]r6\��P��y2�_8hf(�%�ռһY�iy9��a*lD4.\�!�t�U7��3����}A�bo��4�Y��E�F���S_�;����=b��H��5ȥܴg�r&��n�G�j�Hٙ�=ߞ,��PL��in���Qe�g��-��I:��?�q�RƁ�'��v���c�����FV����8
R�� �^�O�m��%�8A��>�pt1@��c.��K-
�h�~X���T
����"��������)�����
)����љ�V_	F�� �~_53�%�<����ަ����5-�d�Ʈx��I1�A�4i-w�*��#l��T�$N|΅[�Dn��!���;2�
M��(/�7�9?�������m1��yz�yڕ�������I�tz�9�Ƶ�SAK?ǯr��ko KJ���d��o�H�v��I��� �l��Zb��	?)5P��.�`�GE��s"�����.&{~a^F䥡�Ι����w�܌% �5��z{^W��?�MZ6!`�5��:���"X��d{#��B]^�sd����<��ڀ���/N������ޢ���+�q-��]�q{���@8|�鴉@@렓�ځ��Lf���%E�0���0���Z�����/.T4�G��X� X.AFp�n���3"� )�X*���cO+o���[OO�:�s�c���z��E��������mDu��^L�H�	Q���պ�dd���@$��������Юr9�t ��� j};�W�3����`��[�$�}>n���ltG5ԕ�|)G?C��0�n����r&��x{J�zSе��zM�*܉?*!��;-^�pe"D����믥�o��NP�2���z:�)c�:�ǂ�Q���b\:&��5�W���o 	�0�7p'�6��;���WCM�6�&����O)~����4q�KP�(R�I"��������-hH+2h��*i������aj�K
-^t���!�J<������ژ{5��r#O��n���R�P�AI1���ޤV����۟_yk8Vrg�#:�C��af� �)= �6��6B7�����	c��c��k��P�R�9p�jC�w���΅ao
���s6�~<	 ��������H&�cX���^n8�NfA,T���E9�R�W{�$@6�V����qq]�t�Ȋ�lP_$͵��Q0�� G�.J�;�n�9�V���Q��%tUB�ǩs� �Ƭ�|���e��h�wƅ��-z� ���o��kl�<k�F�_$Ծ�S71q-1�_�TV;�|sc�a�z��<��K�����b���N�Ű`p�C>���`~�\0aɸ1�+r줆n���y ��Zȡ������'�/��&��Δ�V2&"�֡E*un�h��W��an)&��g�D�A�Q���
vH^�G����MD���=:�n��o����'�/� �dx	+D�U�d���ZB�A��~�8����[��������n}�M��c�{&#��+�����8R>�S.Դ6$!���e�L�z¹\s��j�;%�j)�B��'Ѳ8����PM�\i`+��0:pMu��6�Ҳ�����J��D\�V�U�S��=5A���X��w�ԑ��l�7n�����L"*�Xy=��ߒ<<~�8�ű
5�j�TR<���Yޱ$�7����rR���X����ӥ.+�BtƇ�G������GA��OV���F'S��bA/䂮��4���|A����H�J�ADôш�c�/����F��	<;
q.w4E��{�L�ɻD	�ʛ�Hw=󞒷�y�j2���۾���)��_8�*��&���8��9�E� }:��S��(2�8��W�u���?xۭ�"����e���u&�R$9��IoQe��~�V�!�(.�/9�����f�,� l�m���g�QG ����$K����zΕ���6�Y��YR���BJ����D�d�^�(5�'>)f�x�eٷ>������{Ŷ�L����6�R�{i	Y-b�S�r;�r�P������K��0l���	�I�_K`��#%���ȋ��-w�#�����Z����
�I�	�Zы<��.���:Ee��2�����;$ڴ���TV?�w�^�4C���s�%�t��f��r��J�4���p������s˓�*c�A���_� �����Co����[9�}�t���)ŀt��J��+��F_��W3��b(k1ӏ�KiS��2�X�f�4�� ��y��3�uA���!a��	Xr�֐? �:C�-�/��i*�H"zi�B���u��w�Pc�u���عP�f{>0��R�����_��-E|t�ڿ\Ȼ���EvP�os*^4�׬��N��:���6��@�<��/M��EO�/y(�M�d]X,�9���pd�%�I��CZK=�,��^�i	<'��h��s�O�,���f�wj�`���_�9'v{��Hs#�j�i�Xw��'�\����O�Z ����fu�K�QƃF.t��&DBK�i����hǈ�t]����Y��� ��}�)�ߊ!Tth�de=Wd���'��\
DU�N;�
p9����/�6�Ҳr������-*�� l�0���@suB�~�u26�O�uv*�M5
Ym��l�d�}��1�iV쌗|��^�[AV�[;r#C)�2�n�+"6Ax*Pk����)樹��92N�m�Fe]�,�_S'�B�0��䂾d�����D�b�OB֗C��G:�DB
]��h���ၺB"PH����z��n�,��<�h�V�Y��E��=�!q�����̹�4�-Y+��wK H�˪��ԏ�#��,�k��ǅN�l�ЈG�T�ڮ+�v���>��
�Vn��"�1�O�?����@��Fes�3Y�q�l��31�Sa�\����ۑ����s���G���� ��+�b[j\Y6�����_>����$6Ŵ��}�Zy� ӣTJ�s��Y`@���ʔ�J��i��Y(a�e��H	�;e'@��ŏ�9����n����=�nU��� �$.iK$M�q�(�G���U�������r�g�7X���(%h��=1�\�ቱU��W�NX�g��R�P�Js���r��]���-����Pv�Iq8!K�/V�w�M�B��"}�s�cY��T�!���)��$��^u`���)u A�k��`��
}��"�bml���l��;�LJ��'2F��ZMI�O�:�c��p��~���a-��H�ha9Y��"����������Z��~�Z��\C�g̯�y��L��-c�1��~��Hl�%���å2�4�b,�?"B����C�Zz�C7�0��gypg���V3$َ߲��2�����SdMDJ�1��͘����.{KH�<)v�_4����gO��@��V%�'�s����-�Nc�������l���� ׶%���|����z�O\�3�\a�M���O<$� ��e�<QJ
⽄0��پ�������=�Y��ǋ�=�'�<\�^{�W�jr|�,s;�S��
iT��A�����w>O'�܅�����5�~�;G;?x���0��1`����R,,�d�w���K��p.W�)_+e��r'n��~��Bw�A���񏋧���E�q�y�[�S�DJ�U��|�>w�� �jY��k�tH�P��M�`X.Ȏj��r��^�a^j�x��R�)p�|�~�F�8���'�3�V����>�~��٘> :��w�֓���������j�F�e�@uh�Q1+����HME2(GÎ���Kpnk.Y,w�Ţ=.����c�I~�QY��G�@�U8'l<���H�� ;�⚻{� ��}}[�8���3�z�M���)�f��,��~��x��=h|Zŕ=z;��[��ӻ�E�s[X����O�=�MI�8~*M�Яf�n袍���_�DD�y��%�9��~�|�Qʷ	T�X�!O���,==�`m��-yp9c�W���@* HK�˖���HSG��� R��+�z}�ⷐh�]|�Z^� 4�9E��e��\����B��Ayu���^�hQ����\��6�B��~(��+�
V�=��K��~��[L8J��L�Uco�ɦ�q�"-�)h$*��G +q68P�7�x���5���5�`
�1����a�s� 5�Lr�,�����3�.?H\JGF�5�;4R�#�L�a��J_�#�ۈ�ңwl��$�Xktv�35 *�O�/��Ut�54��%�4L�q��'�ra\�ӗCe��t�{"�o�int���{wg��"K�V&j�c�I�Xj�$�B���[P�`�h�Ea���Q;`�� ��P�R���&
�-����L9�y�W��1V���{0���d�>�(��	����c�#�b*pJ�?�Q�M�&��MF���=+�sl�J�Ś��W��3�Y�7�U9k�U��G��O@R�f3x�x~������Y]�_&����"��µ A��L�\�Zt!*�b]�|�)�^��$����9�Xe�;B���
5�v;��-1�X�3��
3m�9�qdU��AO������BEb��)?r9]5�7�hؤ	k ������"&���@�~�*FC�-9�ua�N�P��&4|�4t��Ƹ�F�ž��)�J�&��,��&�t���^  9��ܥٍ��֖4W]���Ab/�Z����ed̾��-�-ω-B���<��a	aJ����Uj�;��Mc��xtc��q �q�kt�e*Sg�e��{��������|rn�n� �d�	D�V< �R�*m�T�*a�k��ӷ��J��w����t��T�T
�X�%��x�];��yĈF��a�p�cÑ6f˦ܹ���h�������v�7���[RA$��kY�c��pW����<�Az���4~��RDm �]��T=�7�+��n�q!=q�r�7�o�v�9����B�q�?�^��>�����W��@������Y��܀N��!��],�^��z^]3�i�]��{�b���@�����+1�����,8�+Ɵ�v�1�Bl?��$5�r1��4�M]��[<`2|U�Mf爁�no��)b�~GC��Sd��~����o����1�._�l���Ʉx�8�q9lU�����پq��E%^����sSĠ�N߁`���!�wR`����N�e�<�]��e�ZYX�2k6����҂0b�h»á�A��ǲu�^m�l��8hŹ�2kY���f~"�2Կ���e�p(8
�5���i�RƦTGFNU��#�Ҙ�d�(��з"<�I����r�*�Urq�߫�h���Z橏����r��:���6wk=a$f�fY� J�;N����?�y��M���Wxr�-��7��%\s��^͊sY����0n��E��py�<�8�Lʬ4��i74��D�ez�a� yS̈́��#�� ��]���hse�[A*;���K�����_p�C�����P���t���yܒc��1c�O����8첚l��#�\�����C������an��A�s��GI?0�^�Q̊dH3��0XE=�G�jR������`gFw�3GJ���i����!�R���n����."���F b�
ɇ\h"g\#-�z��)w���n�+:��ش�n�7��@�id�	eIc�x{'���b��� /�ٔè����"DdƝ{).{1�'�d{@�A4�d�Xy���5E�٤T��j����oޫ�L�4���[ӴT���jڃ0����]ٮ��=xjpQ�D�x5��u8��U��)�ǂ3<����+�\^�|D	XR����U{��k�zH�@�0�)�[7U R����`�3H��y�"�E6��z/i��#D��d�ڒGbq
7xP[��4�x��G4���h���;.i8 �ySqD\Qy��t)�h�U/CcϪ��H{h���P
�=w H�QئL���^��N�p����K��u��9�Uk��kM�����ü�lJ���~�j�@eh3��MkWx�F�zlϢ�!~�ф��w7����a�#JCqw�i.����b)��b�3���'jN��y�s�������i��b�,�Ooؚ����6�c���Ar��?�����������uD���*��4�-j�"��fV 5�E�!m�s��\�O(9���!A�#�W�uЁ$`<М�x
��x�֥z6sSSh��|r���:�c/��
]"
D��&ˁ�2���i�<��K�Ȟ��fh��#�Z����O,�-k��<�rsU��v�8v�ne���Mj��YN���n�(��-����=�f�<�	�ѡB��e�CՊ��L��i�p����]�9�!�J�^���/y �wH�Q��s��5�x�xj��}�ÿ�gI�x����S&�ģf2��f��Tr�ܪv�L�=��{�W�?�M��jE��wb�Q����w'z�Tk)��� ����9@�W�
<��a�(���.��G��y��zK?�����W(��E(ȍO���>��}��N�m[u�ix�;�͆ր���]$���Y��]³]-���s�)?��	3��Fo�O�1�h��LZ�� ����(С��m'�g%TL���"q�bV����������y5��jjoV���j
I��x'�1��?a
��WD�.�
�<�JK��U��)��6��"���s������ȧK��5�� �1�]���`U�� ��Vx�Ћ�i�Ę/S���W}W����
���('3v)�����@�3!:�_��}q�+}�xI{��Y�K��-������_!��>ꃔc	l8�q��G�A-Mޓ}�BR�l#�Z7�H��Q4w&\�9*��OaM��/��"�c�u�1܄w����C9N={��EG�b��YOT�~�Ej)�j�z��~$��걦9���(w�+.�6�G�8q�򐺃��8B�Xq2zG7�V�i��p��0}ZZx�?T�����-/Y��b5�2�䘧u�Ѳ������*%���7������4��Ĭ�-�00E��Ƈt��v[dX�Z/����߄V~��^VʝJt;/R�w��/}���y`nN��$������Ɣ�7N�@�����REB��QJ��y��0ny�x�'Y�cC`���V:47�'�L��G�I�� ��&�^2�Z�]ȟ�e 
jQ�&��.0 �g�S���е��ZZ��Q�	w�����mZ�g�.�Wg��/Tv�e2,��#@mUZOKT��o��q���e��a�M�u�h<�;�������5�%Ap����H��ꤖ�f]E�| +N`��@{q�cs�f�v�I�총��Ct&����.��&��b2�h)]��z
^0ޭ (�
�dN)�m�ʒ=�a4*��;���J����.x�!%��"�2$�Ȟ��gd��+�3�/1nq*�=^�41����`�ze�k_@?�1?H����T:���u�#��]S��b9V�f�|,?�`�����7��ׄ�n+@"���}��>-_\�>N���_�ܩ�b�FdX�5m�i��������/��Y"�_}F����8:;�e7�~`�!����m�nh�S����-��Id,	�Ҝ ٛFam+Տ( m�R��[���P�f&5�hd�Hm�_�x�~8,gp�F�VCi%�s��CYx]0���c$�;��Ix���8C<���9�7�ja���Ec�}�GKZ����T]�F�݇���Kt��%�Vt����AJMVX��]�3��OR�ZaGD ˁ��:B@>Q��2��J��?oy��ϖ���<��'%� ��pJ�8|�zW���i��z��ÈVJ^�E3�ƻ�ڦ0�U�ֈJ�>�zxl�0n;50F��eo+c�����."����A��yo�S'k�,@�b#<&����Ʀk~��ۨ䍴"��fP��0�P/3{��sՒ#6��g܆Y�R�����ݳ>[:�`�kp̅�(xQVB�m�V"���t��L�gI���o-*=k��[N[q�����p��G�3S�L	�z��T���J	Z�ߚ� \U��5�(�o@�4맢6z����� ���ic*_�A�g�A��_KK`��$��s�^V@�&C�RE�:�� �S��(Tme�L�K�gQ���@(SD��=|vԮv�s �a����>�`��-EKdq:}Y���'>�T��a�����0���|��6���<q��m&nWl�^�w�n��9Ė��F�aO� �,��>��M���?���V��a�f���u­	� ��W�PO4M�NLݦwKԛ;�0"J_{;*�{�o�b������J߈&�M/���p���*LpT!`!t��|W��������⩨�;�*��P��q!�`b��$.�fy�'!R�ˇ�^��{�Ќ@�ʴK��+O��VQM0��աw�Z)����t��+�>�ߎ��Z�*�-VȬz�� ��z��-�2���g��v��[	#ɊK{������ĸ2t����2�8���F�`�ٴ�]��%i֌�UP�狚��ԩ��4�x]\�S�!�0-�w+e���H%��\��"��m{��*�������C	޹�[�x~�&���q�8��;�V.	��-��w�a��4��W%A���0����o��﮳<f
mā�Ƹ�d��'!���%�-�$I(�!3�U������# ����"��k���&dyd��CÝ[���U�W�R$��8!�̒���:#�����/�+����pxI����_0��&
Ku�a�%�C����{��$� ��-��6��܊��~~�/F��1��60���SJ9��D��X��`$#�S���,�7a}S�g��\���Qh-Q�q%PY��u7�����Ȕ`���V�����`��5&c]3&��i�m;[���"�l��a��:r�W�A���`>85�J$�B;2�͌o���?�<A4hn��8z/�Gfw�u8M͹��D�h�#�հ��_�M1r@���Z��4��ˋM6�(�b*E������p����H��ϒi��JV֕77I�=!�zlK���6���{y7�T	��Hb���
�^F>��ޣ�E�����0V���w���3�`~Lo���|�	�];.��]�s�6\ղ���<BN��3���������-4��&����5IK3sr�3R��d �'�mTe�R�6���2���ՋJ�!�R���(�*�H����hjA��`��I�8U�מ�M���*��;Gn�d)#�s#d�D�p�6'�5����W�DӬ%Z�w8�ءѵ�R����g��4+�V�Ӊ��/~D��`���5�7=V��,?��)]'��+�b�P����ޭn3�5�=6�ꪵ!��o�2�@�qđ綬^�����l��/�a����j%�}U���sN�S�W�Ƒ1P s�"ı�wJ��Q����;�.���l�K߉��=�?������/8-�$�M�ibM����>�R�f!dM̌���YJ�ȹ+�
�������z
z���m�����oNk�CW�U�J:�U�zJ��Y���@�\��U���.�l �]0�����Br�L2W5��%��`>�]�Hk�����}�kb�I�=-�Q�R6ɵ��Jh�6��nBA��5��f��<�zLgy�j��@S��5�Zв*�?8 �m�{i�&�`�E}3K!�օ`M�x�Ɉ��ʜ����|�+�/�*�EW��[fN�q�_�kz�D�q�2*�ML�Z�̷�(�B����v�)���XI=��=z�Y�ˍ�����n�w�jeQv�:�b����1ρ�D�n����`^PJCK�m��_� Q�n���?�_.�y��{C�G<��t7�.���f�\M�B �T�m���M�xw�9n���ͳ���:%&8��C ����X�V�H
����]�nˇ6���K��0��aI���U�f�
fS�4��f��@����,��<���.�}��ڒ�N��؈�=�����_^$�k川iI3�G�4eW�J�Q���c[�T���|D��-J~T�a� ��^<x��]�&���Z�5��pß�N��/af����ZM\�CC�+woH��#Xj�q����4F;-���8J]�oi.g�p�hs0=ɵÃ�W��=�~+҉bف��%����۶Vz6�u��)��v�v�_��/�c��б���Piy�;౦S| ^��� �Ѿ�E-`�h��cy�����I�&|�ٚ7���l}�p�W-�M��0M�nnȂ�q7>��/ɇ�Fҧ�L�Cɺe���AӨ�����:cY���+]�Fg�R�Elί.�/�06�6O�|�'.�N�%�)Ef���?��5?�_)����n�+�{WB��-<��Y���۹Z7Y$�aUD�R+&�KD�����2X�	d�@�%�'3�|�i���szG��QXd���� �?e��E�Փ��Yv]Јɩ�7��#�8X���|W�G�F8`�n�J1��8i�
���g@S�7��dG��4�M�]:(��rW*�5�C��� _���{[���5���6�<��"�3��RשR�2��5�e�YY�N[�ݺ���]�ÇҟM�?T�`W �u��ڊ�'|��d�8�ԙ%�9,�M2. �P�Jt*�ڈ��L�3+�c�0u�9��n4Q.���&����QΌXzٿ��l<iSBF�Da�%S��oc5�
fi@6E�C�Eq��M�@�x�X�C��HWK>�VXX�x�ğ:��n[8�S��e]��.�,3��]�� ��1���st�Ȣ9�|'N"�z�뀉;�wT��\q��wp��jBǚ���ϒT�)3m'�z�(�螐�W|�˔�Ο��r]���\=+xs�Q���Q@��&wܦ�ga�MO���G�Q�.����"�|�����������љ�w�56�;����k�r��5��o6<�i�T��|ന�j��hN:w��Z�!� >��f;� <�t:�&:ڙܑB��D�o(>
KqGi.vn��H	�K�c�M�-]����Ӈ&��Ҙ��#
�X#���g�1����� 	w/D4\@ L3�S��k}��qI^�Vʔ�J;ۦ��?K�TK>lЉڭ�Q7�-�f�궪1Z�Cw-��Uޱ�t��hg�V�ja;����ō���N��](��z���3ug��t��x�|� `�t}Y3I؟�ٝ�al��"���٣�� (� ���(u������Gh��������*1!3%�O!+��WV@h_7"/�E��ʼ�#_;���Օ0�������ۇ]�ދ|��20H�kR�:_g�uO�����-�S3O�U��mP�.�L?/A� ӄ�2��<��~��B,�O�$d�f���G��Qr��E^u��P�[�'{�F�`�)�ɔ���a`�������"����Φ0>l'���33ok�ա�5L��&�W�c4�����f��"�H�����G���JN-������)q��/�l��䴻�5���lv
��G>����ij��=�~��*�G��cy�	;��>d}���\}���T�)=,~�H��:XC��7m�7���he�����.��/�����t���֫�H!�(⥐�l�C署7b����ȧ�Lb�xZ�R~r�@��$R}�� =|A�
���5mYUG,�ػ�����O��tL�7�x�k.ȇ�d������ϓu��a_"�5'g1 �=2�_���bP�b5��]��7�3�F��ޜ�2w){]\4d�"�@�O03.�d����d6#��B�[O�"�M�4b>��\$֍C�V�uR1=�����.J�����N��@DdG�ny�����	g}�>�u"������Z�O�E'J�2z�o�7w�+s���y���r�l߆�.r��Ȟ2J�����b.qv�y~���ʐ	g-�:�J���a�a��nl��rRC��G�Q�I~�Z"��|��M���7��
��Q����{#�v���Bw�I)��M��_�i�Pr�C�i�`k���QED�GM�S����X����7h��e��0����`��$�~L�+u�lG�̍[�>¢�2��i�M�\r��M��G�oQ��D=&����_�/+�.�e⪙���6���`SP� ��S�U����pՋv5��f�Y�*"����'ـ��rtߒu��lEBJ$����Ŀ�߾-��ܗN�W�(.�J{)���#�҇N<�&6X#W
�)���(���Z���Z9�����yWq�Y����g�����]��t��_P�H�+���7p�R�x�	������*'j���.��Y���jL�K9ly��v�ք!$�,�	h8�	��_�/����^|Z3{�U6L!�{e�1�J��%������Vz
�>۪�l�K����_cp ��Pf*�����%�;�>ρ�ӕ��S�B�/`��|nx<� )��w����c��V�ޖ� �Jq�Ngh(��?�`o�#Ԙ�	~�wZN����x�`[����C���[���C|2� %�n���Bûs]ʋ���z����{���q�6�q����$y|���s��HϘo�I�2O���U�>����^���>_��8��Z~������>�!�O��{!n'<��H_�c-zؘ�b%J���Wf����r���Z�LV��+��RWo�rɃ�����a7<Ԅv~Vϭ����'*!`5�ǝ�������(~7Z�n��Vp@E�a�ʖ=�[-1�4'0.I�E�Ȫ;��l�<A�N{j�}�[���+�?q��Hޑ����JC^ވ���j��
�q/�D�(��ã���?�&�[5����r��\
�b�DP	a�j��}�����?i4��]��bH�C��.��a���6 ,��1fb�f<��d�G���.�q� ��=��W��x�����,X�~�`�ʪ� ۉ�9��zZZgG�����S�3�pw{%���2[D���҇��*�8�~|O���&A���	�N�����\�s=����P�M`����Ƥ�=�D��pAR�>9f��Ej['�uMn-�+�6���eo�yr"OF��ݙ��B�3`B^������D	�*�(Zt^�N���B��`�}�्1}��������nW<��B�mLMG(�=�ӹ� d)S	���^5�@V�K��?�^;A��-��kF~M�~,�;� L���N�l��h�qU#,7-��ts�n_Jz�p�7̏�)�2�~a`���B]��'�C0��Fg���J-����P�#&[MFn��dk;I�8}��b���$������]�t���������qv���Kߨ�ڗ�%�꧲G���@�����P ����y�o	�,gg���	&�����P�M��(|�=cK��\
�Zx�-�x�լ'������G��$�_��� 5�y��2p^��;��%:�}��k�<���6��654!��Y?��z�ЂD��' ��έ�;.��S]������Q���NH�⒴�҉7Ҙ�5��{ӟ���#��U�r��b���V��@K �N<A��^������ٺ>��M���f[+c�2[�g����M��2��^~�;ib�X��u����OI'�A�����h��2aV ���1�ϊ<�A� W8�6������D�閇��L���lP����EB;&�r�6k�{u����-.�B�ڶЦFQ��+I�þ��1�C�[ԍI�B"�n4�c|�������,�p#�,c��� GCn:5�i��h"��ŬK��=|Cci��9O-ܧd�7�V9|\�[��_]#]`54�<�H[nw-�R*��5�I�y�S�X�a)���2�.4a����GHo'o�6�Io�\�d�r�͍���`�����у���XQ�A�6���fe6�# E��="�l���?i���u�.,.cpP(ְ)�{�>Г,�_'�5����<\a�v���,7���-���v��]cȼ�6ꌴ���\��_PP7w['�*HUŹ�&�[�\��-�my���>�ǋXM4u#T�G|6��Q�ٟ�])̠Q�Oh�Q�;?���&�*�ȅ#f3�L�6��|�h���G%J����Bg��3������~��m�!�"�FAo��R <7����zHÒ�W�:߸\{/L���F7 ���mUy�%�0�x�k+���K�����!�>$���"�J�y��kH�).j����Yw�RGF�ho��J���oj�$\^Ah�]�8F<�q�l��L/f~��#��1iD��,.?�X�e�&/�����_�iR�0�Ro�v5`q<�Rf`IЁ�s_�\��q�*��>]�f�TVfl���Ax�o����Di~>�!���:�x*('�X�\�ޓ���a�����)a�<˱rS�x^&Ve9`{\���]���D �o��Q�m7։]�
�E��5mɨ'qJxSb�u���sH{�-/���>�# �ǈ)f�®Y�rQ ���o����@%�B�y&.�n!�J�J�Ctk�T�(�F7�v@g�uB, t?��䦶Z��)
�eU@�Š[����OG��x�M�UD#�sDּ%̢�F���L���Y��~ug��z�s��{��\�م��տ%aG�p ^�ݡ�+6ۆ3�;�u��0�ˎӦ�Sa屄
|�xUu����R���g^�҄�.��[����-0��ײQ�G�!�Y�띥���8��� ��34o��(R�s{sO��&��$R1 g�KN�5��Ba9|֖����!p;�&�����X��N����J����~
�ᓑu��<���roOU~������7n�)�W#zd7�����vū>��8J�v�3<q��	>��Q"�^Z��Vd�%<!WFՋU��;0Rb]���I}���U:�������n����]�.��	��j�B�cR1E�FqRNk���ܷ��>��a������2�@����d)3�D�:!��۔j�]"uy\_�G6���2�+�%`�>0'�M2�@k��*��_����ܐĊ{�!W��o��E�&m��aY=��ț�M�208w�^12,��]�ihKr�'Z欖v��>9�:� x�dJ��Į8�1�v�)7B�t�y�zyK*��ah�F0�P?7�[��W���$�s������v���k5��G�S����`��h�&�il`��=l��H��C���~,��uۢj�`�5��1#�h�^�g/q�TA�B'��7S�_g��OC� wM�"O(^���kD+t.�/�2��[,t���9ܪ�3�ěP���#fk�f���]�H�V�Cw���.~�J�G��5":� q�hq�`�U6�z/8w:o�<�&i_Q��Nó&� \�%�ci��%�:���L��I//x���\��
�ӶL����N/t�^��f!�t���>2�9[
��D:w�Z�%ї�ag�d
s���zs���dN�%n?ټ�'-�+�4 e�Y�S �ԫ+�鱋yǆ-1L9��ͻAW[�����1p������0!W9��(S�?CnF�xo�*�Q)֛JE����	�a\�V�),�R�0��8��E!��kq��k;/����z�S$�C�77϶7\��W�wr>ЗX#���=%�	c�������a@��CyÌg�������P'�w|?�h3Q�[������$�	3��<�W��;&�[&k�'*y[�*�\O��?�{*rb�m�>P2����R�*o�n�π� P�`�<CsO�8b�� �_PV4�
i�i!����&+b���}��1�Ɋ�_��:�}�I�>>A�H�!����I�r6$��a67na�s��!pa��B喟z��7��
'���1�}��'b��z���;��zk�M�n�u�6��׊����]L��&�w:��ZպoʉbY��SJ�v�q��lz�[��>�}�ܠD���%~�{4L(��|���q1ꇷ��s�*���ٰ?���NA�Gp�J��?�V`���Sp�*YL>t;x�UG�	0Q���ܗ��;�r	�R����^AAj/��^��'ք��&�����b��������`	]:�w���_�yF?,�@��>r���' �L�r�*�p������$e<��c l���x"B�|�{��>������2-��!�I~���hUvC.�����b�k#�R� f�f~m�`Ҟ4h��ӇK����P��Q��<��0���*����wv7�U5�R4�e�C��Y���PPÊ����x��>��O������Q���e\w�
$!U(,1�^�OcL���Fm�u��a���������UA(.�Q���W謣Ka]���`���tF��H��c��9>bO�{����}^z��r�~X�Z*ѡ���a�m��}K�j��3��+4��ѝ]�|\z^�C��=7�tאiF�qr���D�1>���fbR��ߪ�^�"P�|�{��S��쏡��;�v�$�3��M&��U�?~hk3 ��5�ޘ${�D1홖�|!\��}�3^5�a�5'Q1�2�Ǣ��46�@b!��X�/x9pK�,�r3���j�ˁ!'2xlK�Q��D��C�O���,~&7R�� Ru��1�	�_D�&;��_
Ɲ~��nʘ�$,ңHn����m1I�?ѳ�{��Uu#�g1U�S��ݘ�ȹ= 	� y����пk)������;�G+\���������K1�J1�1uz҄��řYԸ?��o�7�X��.BX���e���� ��;J��k{%ɑ��~���W��+V?@~:Yi�JE�k$���B����"� �b1��<�8�G��d��`<PG�O�,�AjM���n����ܧF	V_� ���B����3#�L�Z]��:����N�
8k��{i��rE����^�D�)?��M>����)r0��\���o��A�<��Rț�{��N[DY�K�m	j�&��ɓa\�s�r��
�*�nCA2N�fh��6���/���NCDŽ���G����Ѥ[��>��R����7�x�^��͢�b(%���`5�^�$�p]*�LL����o�s %��VR�� �n��ڕ�\�	�nxiڠ���>����Է4&���4�#\+�"}X�%�K���N�������/p�f_<�B�h�-ӯ���'F�W����uË���t����o�"�6~�V��\��qP��ۥ�~w�G��� ��j2�𜖁��$�T���˖��/�L�h�$Y�/���t
����2>滲��m��J]Ʉ��?�����8��-!v�o�[��L^T����^=s��f���&���>����S�E��0kh%H|����������Ԕ�[�({����4����n� �Q7�e@$���8W�C�0��!��D�D�h��Cn~X�w0��Ğ c����GcE.�v��!Q��E������z&��vT��~I<}K��P�@�'��L����k�@�\�`5������e9�r$��}nV�I�,I��$�d���|@�/���"0]��(D`�E�?a?��6��U�<�2��c}mu�d��e瞹H8��͡��8�*%�	X��xi��? K�c�ٍ�b-[������'��B{q6_�Cݱh�� )����䜃�c+UW6�*����+��:G�F<!Zv�Z�;�FI%o9Z�qB3��2(�ޣ�"T z�����_��,A\ș��k� �f�1YDE�DC��xХ���	�30gLYn�����õjB��Y����4bl��k��aݕ��1�o�9��0�����9Q�)��؅��\��Q�����(�1�M�&�k�L\~��z�X�<��k?ܔ�кV�wxR�ͼi/N�{V�[+��ï���%=�d�	�n�4�T$�f.��������E�>459�d���q��Y�����)��Gr�&x��L?[?iX�/`���܉�'t
�E�7�o.�=����M�%^�fS>�N�B��y�e��]	�e^t}�ľ�x'о=XJs  W@o�`�nu�J���뢻Vc���gjP j�$���a��
��S������ղ�<�r_º�m���6L�a�0����γ=��n�bx�g���X�ܢJa2U�ȕ]�6m,c�UHc�y[d;�6�]|����wG�ԡ��`�L頬겯[��ݦ�������B)e܎�j�bѼ�[HTzP>9>�s�U����S�H�����M��N׵w�-���\a�)*]N���� ���R��ڳo#�k���o
�IpT �Z�m�IX^\j�j�A{ڛ�#�O�-����i��vԺv��*g�y�Q�Օ��쾶�ܻz5ŭs��D{r˸���z)�lS����eK�PGw堂a�J�?��0��*�W�@:�$*��`�;��!�[��l��cTbQ���6Rx��}�Rb�]ݙ��BF�)�g�&����$�r������O��'$�����7&�����[=�h,�D�UeaH�t#l���O�̟a�<�� O�y�*� {Zs�}���:'���M��C�F�M�C�}�	��y�kz���!6ReK��B���!(E��q3� �p�.or�����(xXn��Q\9*'%Բ���Ǎ3�ǸGV�Z\#j��}�HD�?b�Vy~7�P��D,Ny8+$��e�dV�����fYO^����7hH��J*��py���8�Q8O&��ps�1��?<8=��<�a�����7�0`EF&�ͦݦ1�����R���� ~������	��ШC�����s0��5��*)��ч.G��\�(�Oo<dG��)V��y�*2Ӣ���D��L�}�+����$WvEl3~���	"m72��[�(�~	D�v��:-��,f!_�v�mB�'�Ab���i�%���n}����E��3�6�nFw�m��lYڡ-=w$r��Z�
 Tm�'�g�H9��K1�0���!x?^���"�ƍ��{R�*�s}QBԍc����w`�p�G�q��޵]��P;�գb��-~��U����尙S$�<j����%WVg��#�� ��-�JkKN;��8�$�#������s���r����-��"9p�Dcf�T�;H�����R0!�g���d8S�=I�c�%�rlW�>��=Â�P�cK3j��Ħt�O��l)��*�͚�1��D1+*cg�bU#�e<ܢ��o�w/��;"B;-�)4 �N��?t�����?x*D� ꊫ56a�W����T�[����8��o�2�R��~bv��R�x ����������8	�"B9'�7̮w?46n���������,K7�RH�D��V�y*�F�#$fj�1]fI��ٲ��z{J,2&�q~%8O�Ag;Fm�+�2���6�H�u�E^��g�X����r�	R����0WZ_�&���<0귃��)��%�y�̟�p��<�"�=5�ĕ�!�pǟ /1x�2逦a�n��_�dPs x	S��=��iRz�8P�=0p]�+Qz�]_�u0�
� �$J�*���QwC�U�ћV��B
މ]~b{����Ճ�%�.�����'�(�0��J�
o�n���~�s9��˂}�<��b�dI��K/{�7���9]Z���e�z��WD�=rk�)�#��LZ-=�Nf�.�'[�̥f����h�u�J*I����Ai��܍�Z�:i�S���O/�b�V�Ͷ��2���6�2�+��@$66�(\s�2�Ԭz���HB��%��]j���8��i{���-]߱��Կ5�S��&,�.)���L,�f�·ˢ���7��1�y(>��0��w���W���4w6^�qq-^�!�2gO�dy��&Y����[�̔W���\��G����ߖ�y���'9M��G7Vě�TWcs��2 ��񃂯m���{��?1^�>��z6�\�W���݅㊭w!+`���s�f���=��gb#�k�}��;�~Q���d��W��ѠF�Sa8snK�
v��i�s��7�bF��ٖ�]�.������Hens-E<�p�҂�k&r�� F�\�՘XY!qTK��s���4�5"n�G�5S_o��9�(����g��S�
�8�~F�[���q�U��g0�*C����Ce#U�*��n�!q����;K� �B���ɷ{6�/�@�?��9OjH[)�N�b�<��M�S�����t�	`����w�"=�� 4f�P%K�hG�:xd��j�����GO�׺�}ߝ�%�^�����5������["jɄ�r�&�$��F�kڥ�]BO�[D�xo�֘�L������ �$�IH�e8\���A?���
���ԭ�ܵd�t
��t0��E+��2E� ��)�[ha�\Mޑ�Nr�+���p����2�M��Ғ�8}
���)����F^%���2�iZ��a����   !5,���И��~ا^ĕޗH�����q� >E�X?��<݆�M�RL�A��8�>G�RwJ�s��:���z�uikB��[0���s[� G�V�G�P�.5}!~�}�q ���`d��E�����ǥ�*Ǧ�]w��Z�Y����˛U���<�dT�On	���&+��!#���<� ����Ư"�� DL��!/zlt'5c�S�b%�����PWr/�m�1�X���G�)��t6eG-��o�Y�,����D��%��""7���_?�� ^����u�e�ŋ�T���zx[�����a+�8�K�\m�I��Sw��YTܗ�"���WQ��n؂�eM�JJ�5��=�Ǌ4L;4+XzsF%��:��򎩞���%�A� ���h�h�F�8�-�n��Ǒ)Qb�����si47qd�nH'�}-Ρ��k(���UA����m*}/T�)��
�|�fpxwE�6�4�������x��N�G�H>Ϗ�j���U'"�s�Z���@��|/8S�ob�[:5ڹ33&�[:s#��A��rh��sUn#,R�������~��e?�Pd��{ ��݁8D�&�kӖ�4�T>�D{�6k��̳���;�kc-Q5�40�"sc>�>wi�]QP-�㩯�oi�h�;5���ڌ[L��y�:�(�0a�l	
16������4��KJS�����O�^��Hb��B��SRKy8&|8��K3�L�����r*��8n�$O�����ݼ��A��v ICR�)�UJ�x�*%�&[�:,@�;ݒh��+��p�d=Ʃ`��8Hb�h�� -k�5?��s)�]�n4D�BB�hڵ��t�b�r��X5���>�U��!��ch��V���þ�)'/����\�fa����%f��^�&.�G��h���@�X�>�[�;"�ޣ
��{L��{�s;5�l���_!U��`yONt9n�-\n@40�6��`>~+��=8L���2�~X��e]�$�P#���W7�ڕg��H/bA�޼b�C�i�N�g�F�����C:�� �ԕHeP����갗R$�8��~\����P���C5������j!R���~tۥ�Δ"t,�˂�|���7[������g7a�:d[�jcs�z
�(�m�ؓ�5��-rQ�SC�􉆠?�ؓ���
fa=3��̠}��Y"a�i����S\X� ��7��M7:�.�����U�ژ6���0���σ�/��]��_�����;B�*-q����v���۹���R����7i���I2�	nGhiڐ��5^����݂��^<�j~���ޟ��\Gv�۩M��|����rrpM^JmU/۫����ط�]쎦J���W��g�b����&]�ޅ���rU�����6p�I0�<��n�3T+���+�{�g���:Z��m��T��0�[�S�?Z����:�=h:iο�Ic.�I����4���+��
�͗yr3�O9��|�Wպh��1P'�3i�Uu�#Z@�y�f�]��������yr��(y�x�Ny	Z�C^z�+�%\*�KcC�8�߼�G�VC:xՓ�o6�װ�;���_���I�_���6?82�J���|ڊ�n:A.<�c�j(��=n-�.�a�G��4O�40��KA��a�*Ș��]VІ�1�wQ�ھ�0�b�͗������D�l�ЦVW��,Cє]�Y���ɚ}h��aO%�,�U�-�����ݮ�S�7��U�I���x�6��iW��l%%��*83��Y�J�@�$��4>F�DO!�� �l_*��uK��y��18$�ņ������;�t�ݡE]���2uS�v�,!��cƕ
֮ON��_�D{�ک &2p��5�ł[�ol�� -���9�M����a)t�z��t~�A�$��VJ������ Ī�2�j����Ǩ� �Bp�]�Q�1��d��]�5���j���oZA��g@���V������q��rt��SX^�5����9��休	����&{���beIkF���SEs�� �%��Ȑ`O��N�"��aI��Aѽ�Bb�u0��F��1�M� z?��Gz�}��n�РP\�d���^E��p��<��[A�r��-��k.��_��Ӣ����T�� =�.聾�O�,XB�ncx��F.�;�Y� �^��8S�+� v+�!�s|�w�����,t)]=�˶�5��E�#���ƍ�?!w_��Z�L��d?� �7t���7R�2�0'?i��P8��#x�^�o�H7A��$�� 2Z`s�?"�� Y��톙�BUoHSU[zjVIb9د�1���\���#8sT�v�'�$�`�����.���;�|Y�H�z]|�N$���Sc,��d��HF�8KOB-����,%���a,=]&!��M�G�gU~������Xw�l���i���8?v�T�p5�C�^f?t��|Q�e�F@Y���� ~��X�
xΒ\͌3������^�ң�Q��:p�,N�!s�5X�%B�	娶��3����`{�|�5QLm*����Smv�:�i����2��[l��&���f�=vw�_I͒gj�m��n+?�!� �YM��B��OrW�I�����(���Xѽ��C�g�K�/��Erҿ3|�u,K�@w�Ewv����ޞI���Y���Үp0Y����n�=Ij�8t��`�݂��A�K���J�pH=�<�Iףa��o�{M����D�02���+`Xi�w�i�wB�\&�HE~Yڗ����`�l%�M���b����	�����"@w<�L���Kԭo3�� �w����w)	�[^�Y���^z�/8{0�9J�������_��b�4y�x� b_��Kv��N�(]u��I�M�H��VpbS�&���yc�6�x��� ����k�JHL����1���a���X
��s��F�)�u��Q�T���~�ﳬ���zlw�: �{��dyen�/mNS�<���Lg��Z��Y�X�w Cx��1,<�N��R<�ԹN��� 4.&jC�n����d!>�Q�/�����)�2O���6o���I=�G�G_X���t��΢4��ʺ�+.L������Y��'��<\|cd؈䯬��g�~7�H[Me���M���~ �Wf~��g�bd��OxB�����y��!R���@r�C��eb���\�rۂ������P��vN��eɅg��CMI]kVD7�]�)��Ʈ�����1ץMՇ�ɰ����Fl���-��Є�~r*�J'��t67�*���y��M�VQ����{��	V;�Z��zHʃ���@�ҜÇ���be���+[~�J��w^�<�U�ҳ��n�q��;g��N#E�&����>\�6��k�P���[��m������5\$����D�DE�������D[��Б�r��
&��LU4�!9���.a�^�&��]L�K[5�[?yҎa[_�~���T&gӀ_�ҿ۩q���"��D굑�*��6���Ȥ�:��ޅl����/���9���9 M�O~���=� �x:�� 8QK����d�[�q�B��r�����б:
ܼ$�v9^�/��̚�Ҁ��Jĉj�lo���/�����Tߚ��^�р�(ia�x���]�ǆ����l��;	�9���r��a.r`bۃN���K�V+�� �(l���px"�*V �f:� �b��^�a2�/�U�Z�Z�pn�Cs�\82Wg�9�9���C'z,�*�j��,*\�o�9N쏼ߜ��*i"ĸ�d�TDIl�h���A���f�{F�Z�\N��@��~�~(Ӫ���#����=�"x�f�^T�D#M~Ö~n]�F̴�����b]r�����`^fke@���[̂F�:�>���k+9ګ7�8Z��O�;��~�ҽF��5�WjT̯���D#�z� (H=����}�ۼZ���~J�!sj��xRV��`�u?e��
�h��}��}^�mZ�'����CC�������J�X ��xp�aR�YZ���FS@�	��ΐ�S"��%z�}��Rsy׿�f\YO(�0�1��)̰��^`����$��Jm(�ke#b�W*[_eb�@��(8��,�On��(e�mP�,�c
!�[��?,'_=�\�,{�,U[��	�1(RW��f���«}+�hw��0#�U�}���Hm�9@ΖC�q|�g��+��j��r�@��^���-��ȅ���k��GΪb�C�H�eI4%��.���9W-�\�p�B��k��x5/��[����,�1�6�Ɨ�&�*ׄ��lE�0m�'���I̷���^�!.�˯c'��(���G����r��$�iT����r'��K�ipB<si�U��F���$X`���{T��ڙ����'Y�ͲlYD7t��|���U�����b�w�жIIđT�O~�5�M����?�q8D�F�w^�+Y `�� ��$�?������y�&^ԫ�|]��v�֮�۽�F���*^��g2BR����6�>y[w��feB�.�Ԁ�ʆDi���|Ђ����!?��7�-C;f�������O�(P������YCB��n}���z��JT"�U�F�n�6t���;�%G�yԪ�LA�si��_�G>f5F0ޤ�Uш���R�V�}�*kgeD_��Ɓ�:et'ӭ}��|��n�.��(�D�7"Lޮ�[?�z���]�1���~=j�:�n��#�,Ƹ����W������;"� �;R&�r�9��yn�������ɫh_�[���7^����N�.YO�1���fBhQ󫦃f�?���X(w�Q�C�5�f��͞C��%����b�-e1������;�2�=����]�w���yi�@�w���0�FGG@M����3<�z7\808N�����s�U�sX�س*�'�UG!������*���sU�}�rW������7o��'���p.n �t���Μz��:�nU�N��R�!$p �ܮʺa8r�?�ŇD4�g�6�������YGQ�o�O�0��<қ���O����T1"�
^i\��w������G,�>���
Gxy��Y_�!���P�w�Z��ue���nX��I��7����1����Я�Ѐny,j�c1Bt+�{ķW[fItWʍ����nʸ[D�*�W��q��6ϑ�M,g]�/ۧ]YyClL����M�'��6�Y�6a$"�TpN�f��im�Θ5��0_G��t�]�����e���$N^j���%�w+�hcg�]�����@7����:��J�VYS�1��Ȥi�79/�ؚ�KxB\�ֆC��\�����|��IN�ɦ�s5��©�&3D�8k�̬��#���_�E�l��o�T3�Կ�'��\AR��\�kj��y�9I���ᝐܻ �B�����!��=b���8�fK�J���qV�B�s=���@5l.iRM��c��#�3�p!�9N����˰���N���jlu�5���+��c�\А�ûr@�k]�&�7Ղ!!�������}���x�n����e��I"�q�$T��b�"�v5���1�"���8��c�d�hhh�Ӈ�;�AU�-Q�T�����O�&��^�-���.�.\��K`C�so�˞{'���R���n�BD�@B��+���~���(����U�)^ɤ�l eA���N���Nb���1W�Le[���P2��L��B>�}��.�bNG)������� x�;�յd�0퉆�ɹPz(�D�{7�FV+�T�f}��p�&J�A(O�~����fE�ʏt�5�';��N$����u$VU��ˈn��I �m���R�B��s<&Zێ�d5+ٮ��f_���JF��qKq��o9��z�c��o|�OS�G�OR���)�ee�#�쿮0��b�ě���O�AA�[W	m�������$O�&[Wd򨿄"�p�$\��!>W�����Q������E+�-v?y"������4��6�&>��؀�
`%�mW�J���F��>�챽����ӥ1.w���k~�k�A\��$�TXD85��2�~��]�v�6�&P`X�}��	� �B�ns4��!��Xˮf��ߟ���SyJ�-�Q8i�İ��$*�	�~���5����6�^�,Nt�ɢ����[+�[&��,��No��#9tw���N<�
5�k8Ij�g%� )#-آ�[g3?�.ߦ �
Ӻ�u�X����(�3?Pꧧ-�/j�4���mr@�ޓK����E���LC��#��+;��՞Qg�W���g��o\�Kj�GS�ݳW���C�k����W��Y�� ��	>�"k^; �^� F������bRQ���~?�iu�^@9):�X��1���2X�)][*_<1Os�(z��}I����y�)��c��-#��^(r�8.�pR���Y��"�ZNt��u$q�xIIP�:5�N�P}��b��k�^�8�Ms���]"�_9�c<SH=mX�^�2TLP
��[	%(�3���i��}_��opL8�����N2�j6#�wNvRL��F�ù
�2-�^	c ���E'8w\����#��$����uD��~��a�$�E0�#|_��M�,`�I@=����9-,��'�!.o�v���n���#E��t��R=ќϧ�L4i��vJh�e�[�9FX��H�.��f�d��]e�����d/��_f=�γӑ���E����f3�la00�|�9ٓ����
rZ�����la� ���<q}[���3����ݗP��W�����#\�?�O���<��lD�J��ˏI��͵���w��BL�"��~����ͩ~��_�8��sl��|�`�&B;[r	E�'_w/�������<v6qEb�oE�o��3O�i��P(Y�).Mb�n�Y�[l
�؃�&z��1��>��P���B�7�(�Ynt�)<�/��ȏC,�٧�5��z(��m��;
`z�Al^���mUP��{�+2޴Q�_,@Vx(�Ǽ/�Dv���E\�S�$IO�K3̊���0b�R����V�lY�;F�i��%�4q-L�ԉ�L��^��G�J�zq������<��qm m9t�x/��@���a,f�g��q% �7�8>��$�7�ܲ�����-Y���C��*m%�X��,	����#kK;�^Ά�&wcx�`*O#fj�H��{i�(�i���{? 3���8
|տ�El�@����C5i˃��lU`��G[���Kz��Ҥ����){G�s#}�ԑ]Y��oD(�W���P`��=Z� w�(���+�m��������m�<�OCU�b���W�k
��+�;p#E�Ϭ�1����MO�na]w��@�����_�4�.2�8nJ ����6Kt �I%od���78W�xI�J7'�PV�J�G��v�䁅w&D��Y�uƃ�h(� w/Cp��l;�ņ\~�{�B�]�y��/ƌH\�c���?R/�
E���|/lDm.�sK� ��dĜ�7�F$�u5���?M��<ۮ��.���l+2�1t�o�D]���Ru��"��h�'���̲ \�uuPl4�R�ҽ�0� #���t�_���=��9��)���dˍ�cn�(��8AB(&��]w�+��3��ը)x�W��R�\Fxue�k0p%��n��[�5���s'�;R�lv+�A�gx��A'��7�L����Xy�����&r�i��������Q{3��?��\�mb���|Ԋ����2�?�u�p�TaH�It���;ڂ�Ǖ���~��l5'��m}f��v�j��(�Hnx>��m3&�܏;YSm�j@R��Ɣ����t���w�I�Y'y]���a�]���� u�Qhh�c��+�6���̙�7,v�����X6�*c
W��Kԥkc$+Fe)���Q���#��t����Z���< 
�%{>@�X��ly�ƧY��jm���K�"	)"�.F�('��~��D�B�}♒O�Ǝ��n(c�>��8p�	��V��D��|�_��7(*�U�F�� �e��������H��suw��k뭠��32(�V��s�D�����p��!77az�������f�A��&W�3��ܥ�H��ΡuP�]>�������k��/�"2������0�D~~����ܺ���x��%''����FB��;��F�>��C��5c�V�C2�ǳ�
�5V��
tDE�w��LK�.�7�n(a�ᡪ�� �,�A���F~5��� o@�� S��{�r���:?���Ѩ���S��2���W�~UeӕJVUL5��z8�[2aU;�H��r�]�"��������>�ʹ�o %�^̶�e���ِ �V�l�D�
���ٓ��l
�-'��{2���T\ך�} �%��*�6��9���s����O��9!������j��p~�V ����^�7�sx��w(TG����H��c���!{��!���dZ?Cf�h&����\p
"�D�i���kT����J�H4�e�B��~�j��{a2��s X�Wu�ht)��t<��q�\N±4�e�']ED���\���Ը��$��^�s�	nó�f�/��-�Л�r�5������2d;
	ª��~�A���!�o�#YHr�T�w�`y�G��r�"ʔ��a����Z�����l��t�޽Ǿ�Z:W9K��DU�1��W
����H��\������I�II���Y*��?kq��o��UF�u ���Y�#o���X͋̽8#���i��ܮW"���]8I-L��s��8_���W�+i8�:pL�y��Ŗqƽ��&~�d�}��G��5J����fy����M���"a+R<�B6{#y4��]������L�����[�fɜZ�䔞�ד�#�5�mB�tu/E�A�Lf9��1�J5�<#-`G�	���pQ�ƃ��O{�G'�=����Cb��*�?��Я4�ڱ�ͥP�׀��4?�IQb�V3�-Z|o��9X�Ȫ�b�.jZ��*ѐL=�b=�p�^iQ[��VK��fǤ�������KC]���Ms<SԨ0.�G܂x��V(�����3GIY��v�F��I���� 6��md�Fw��H���[

!/*��A�%/�a�����0貐?T��<ԩ�����5$�M�ʿ"8�M샾��*�5��H��,�b�5�F[���f���`�gܠ��mEo�S?��e�œ̛��y�L�q�\��!Q�o��lWV�����0��-�L�he��U8��ʎU��n�П8%,�?��2@ͦ�|@B��Ep(^��מ?=Qݑ5�"�b5|�C��AbLL
U9d������;c��ʳ���,���.��Z������O!��8sg�/p��w�obL�*30�j#��bU<�o [L����J����l{�����V_q0 �) �u����0���)��-m���~��3s�΋Z�"�#��q����;����N0"X��ŦQ/�6S���*�R�h�Ե
�qq`��:�Lܮ��3���rv��j���ظh�����#1.{����M��S�w&��yض�+��g�	�n������]�P���2O�*�)���S�7A~����_�=PmX��9;�%QB���T�"Q�}��<sƐ���^�}�<>�j-M�^DC��$I��X:2���ag��(}G���`�`���]v���>�+��r������E��.1v�y�js.�^}�88H�v��i;Dc��6�~F�g�@�nт6��T��"��Ld4q>�A_j!|p>���-~�����xp4��&�Ȣ�q�p	����h�P*�X�@�[�W�U�(M���k�)���%7�I�x������+��O`O��s\�\ր�.l;��i*Ǳ\�
{�!��Y����(M�/6�����rK2��dd�>���ЀN"��-ވ"w.�!Cb���A��96F;2���.~��_)�0�x��m����*�� �3��u�;TJ(�^�#�Y�C���Y�L}�A3�C�=JaW�8D�HR-I���N���jV�����'�R*Eʓy^JCb�mW��UX愆VB�G�k�
����uZN5�!��C��oX[>�!E�;_>8�`7ǖ�Y���~�J�h���>Ŀ�Z�+=�P/V�m��Zk^�˅���	��ǐ%���}�rywcգz��7�#��F #���DZ�4��v�]���D>��x�eM�����8�N|h���|0I��`���&r����vcL��fq�s��
�VjV�5;��ƛ%��:C>���zGJ-����#�4�UPNc��m��t�P���rr��"2��k��s����Q/
�&�3��HK����g�e��/RS���3-u3��^ï�Z���E����Y@��ޙb@ag�����H'��&�#���.:b9z�9g 	�����呫�&��a����@�;��΁P���2v�������&>�N)U�
�7^3tv�� u��S����Jȗ�d}�vY0�Oc���>J6�3x,��B~�i���k�>"Ř�&��#'.a&A��E�"�R!`� 1��9x�=VIv0���ZL�I��-�3��؀;�m�8a���;�}K�+bk����ն�L�}1S�Z����
�r'�v-
�=�fԩR@�%��ڗ��:�m|j��2�� �b�����2�t�A�_W;ҰzS�>kZj��M SkAQ E�����A^���."td��"U�c�����C��X������9�ކ��s�L�����ĥr-�<՗ٸ�pE7T}� �&Q�n��g<\RQ+�c��ޗ��gk�=�jʋ�7��H���#���ׯh8�3��),��5lP�SS�ϗ��dV�߰�����u��Q3��Wg<cL9���l_3�&�.ԕ�:Q���,3�V�7����rq��{aN,���
��VX�5�Q��r�Zn�����޵�]| ���${v|a��(���i`��m��u����Z8!���x�Un��EIa�j��Ud<�U�a8��F�ZH�^�hmx)�������$�uŲ�zE�C�G�c���j��Ⱥ�W���h]�1�
�+�|k@�M����}x��:��=���a���e�(y�<l'`�ԜP*��
�@�yx�)%�
珓#\}�?��]
��S֐����� 7�KR^�= o»M� ��� [�]6Tt��z�9\���>���c��j�WqޢpV��w>Z���s@�Ot������so����B���HTTY�h�:bv@�i-Do<�|��<-)tP�%9����ep���B
���s׾�.�N��*���:��j˝�h��syK.��oC`���=��/5���eD�L(q:9�c9?Lf�l�"=^�Ԡe��S��,R��9��	�Ao8#�TU�9Z'ӆ��y|�T!{�ē
�����8�P���swe.�=[�#��{��hT��`��JR���E[�M:�>�� ia�]B"���(`����� ��Ʉ��q�v�,�ʠ�@X��������`b�n�JX�A ����@a;�w;5sa��5œ����'���y�Ip��[����\⳶�JG���9���99��P��řn�}��X%�[��ԭXOyj].�����N<�Ҷt@>����&7ש嬎խ.D��
w�ڝ�'���L�ǉ�}a->���<��̴�ȚUҺ��xJę6 N2�	CC,�5�*�y�[ag�}_,�4x�+��y�g ���/�1����3�e�@?��P��s���1	�X��5��10���ݘ;�ჩ_]�rf�u���\T��m�D4dU'r��zM\e����"ʓ����Ps�����|��zn85o���[D�5X��8�w��,`�ɣ[$���ٕ��Ojfd��<Y'4W��x�O�ϧk+��$�Z^��!��b�ĳ�c��}´e�qͤ�r����(��� Ҫ�ȁ|j��@	�
@�O%���Q&S䏦t��+�2�Q8�]����D?��+������<?��4'>�Gkٗ�ܚ��1f7�\#K�+@k�"��_{T�j�/ٶ��S�~��&���)$i���'
�x_�3�t{���v��Nb����c5$�}��Z�%�������i��*���/>��Q@�cO� aR��6�Pvî߱ͻ��*M���*�d�
��N�Z��j��k<��J�շ~�}�	�m��rd�����;S������|�{�B�EE�h���q��9,Ζ�����=-�<�u��y���Qnr�[y2Pi�zi�2M��ᰟt�6�0����f�
��I��D�~�Vh:���
�`)4
0��[}��hh'��Q�W����J�ʃ�;B?d��C�D(O��6(�5c 2bƅ��Y��6=^�2���!c��D�m��_C@k��W�k��p��煄�����2��|���V��Qi�Ȗ^	���w���;�N�����e�vSH���X:�'y���DfJ�*�:��t��.����";��(�uٳ���T�s|�8�w]U��UC��&^����a����Ф��,�~����,!VPi0�uJ�"M;C�ik���2]�*謘E�	�檱�*}��\Y�q�-߯E�\��V!s��<�Ý�	�7ભ���߁,*L�Z�v�M�,lLߝ�hvӳ9���S	�0o��W���j' ��l��P��9R?"�=E�v�U� mO��t ����^WBKK���S���Bq��6�襐7�ȫ�j�]y�2աQmb���K��żFʀ�ë�U�7l~�5�i�u�Vנx�?�2/GF��D��%��#�l�V���e�=�2�/�y�Ce�Wl.����뒩=�� ��\?	�K+��}���ǫ�TY��8�%l#�l_w���/8���~sBN�'�fr��eȨ�+W�I�簿;��z�1���U�u�©��h�
C	8Xi��2�fOYtq�Dڍ��8eԉ���Qw�y߀����1A��i����50���Ĭ��i.
4����b��	*�|7"XI
G�q=�����c���},�ԛ�Nv�9���� ��A��An�h�m�{�/�qait�t$�\1��� j���AQ*D�st1z�����~^5�!Tt�͉j�2kl�5u晖��fij�u5�<�����V�ܜ��&c����*z�09�`�#��b��?`���4�&�=����QWݪ��Rb�c��o����>��}\a�8.�{0qjN�Z�Yp�M~*�wR�CS�
��L�;
fM)�x]����5R=�3��V�/\
֞�n�*R�>��d�ɦ���2�aU~�=9�G�����7���8�xs��l�ף�س��!���|�J��Q��WҟM�G�<}�c��`v�s��!�\�H���4)ؚn�V��'�s��N�#�� �!*�H&����WN{���j���L��D����!&�D1ԗx��tf�.�6���e����94�O�|�T`)v�{g^t-��xeկ6�u^T�U6m��׏Tt��c�m�f�T��|%r�+�,w�l7��m$z�sQ��������.��U��c{�Xf�O*��,�Σ��R����gυ��U���ܼ06Y"@@�+nx0>�7?�N�K#�5Oe=��g�L���ҧ�AT~��-+���^y��J��Qn'�y�/5���t|�7*��v��P��oZ�WN|x�<mI-�׷���٩@�Y7�ΡG��R�CO��$k�M���(oG_@��鵯�5�D���I�ƾ�E�`�=��O����h�i!��G�(jO�WP�(1�5�z�8,
T��`�X�ʂN����`���Ź��������'��L�C�j�8�n�2g�4�.@��Y�Aq��X�{ud.NxW��4���@~JJ�.��"G-��j�ƛ�=�%Ա%7��Ǫl�Ҡ	��.��+��� �;P��[E'rz-5��{B����>k�GD+O�u����2�t�^F�s�(��1x°�z���7�L�W�\�O��D1�J�w�m���mN"X��d�$T?��Py�ViJ�Yڇ|vcj�]�̦��Wo�_��`
��6ӡ,B��X�7:�����se�ĉ��I��?�&���p ����]���>\����ե���Q�������D�Oj`���Hd�n�{Y��>n���N���@�TI
B���:=�ɜ�`o!4r)8s�P�&�o��B�9I����0��c�>ZGti�3�T�!,�s&4��C\�{x3\e� ����'�w.3����j[M�ű������Ӻ �^����`���~��j{�ե9+u��E�4?D'������jZ�q�x��U���0&_Ҡ��[s�'�ՙsj'9F�S4�i렃H���r��H�w�<�p;��؀�z恪�L.��_Ow�O����!J��&�@Q�<tm��(���#9*t�A,�f:�aӶ!ܚ�K���1�����(i�@����PlB���s��#|�9sZ��i�v���0��j��v0p�X�9W��2�ݱ��D���x?����h�vbZ��-�D,/1?�8`wi�PT��[X�N�a���4��@zkB�2���JN����u��$�}�!B9�1�jSE	q�&�t��yc�nwQ�t4���"+!���gC����_����T�1�J|X+�z����:ԍ���3
b�K��T�B��CK���Z�[��'��E�S�'�t�xN�5
���/�5wT
�i��d4K�֮ݣ�6��iݷF���q%�%�Eº�9E7����Jf��Y�kb��c3�W�**��|���m�;��"g�	�<���h4�����{��4`�fr�\Yi����\H�h"5��X��z�!p��Yn�]��d�\:�߀��/�.�#�g�wr�N�f(��x���#E����M���K�`�(�u��#����^06h�H�ҹ<��"
��]Cŝ����,V�7�ϥ*k���cd7�}p¡nȒ�"�
��X�����(�e$��9x�hO�J
C��m�6% �_Z�{K]�?"�f_e�؋�d؃�t;,��eҥ�C���f¬�/9k,q�^���e����-�Qs�[���pb�d��6x�Y]e�� '�g5A��L;��b�-{���b�y8�m�}y��v�g��}����F��T��	NU�I�«Y>8��!L(n+5[�ߗ���
D�L�e(1��v��Oh�J�AE��I�c�|q,B��vR������Cx�}�*1Y:c��P����eo�$�l���c�3y������h�B�l���+Rq���-0��d��Z�R���u���6������(=Fd��,���:W�H;�gC���ĺ��'N��P�Ix�!q����	��_|���ͤi# BY�>��ɘ�m�{�ҥM5�s�e�P���)�e6S@=��&��R����Ŧ�1��R~h<=�޹�� �K�)��r�c&��(��֝�26�o�/E���T˹K�]�B
�b~��.u���v���)��a�eX��͵I˶t12�̋D�-�C�����4.W9�L4�Ȥ��0��Q�6P������ʫ[�e+��]G�`�шWL��L��S�3�G�ꎨ��,��1-M��O��37�5[JV2��<wz>���.ן*�d��H]��ﾼ)�	�k��JS #3MV[_���$ͼ�?�����+�9��(;Z�:5�y��b����*��"��^�-��'����)��x��� ������
�������ڼ�¸r<u�v�L�����e2�q<C���w<���ҕŰ@r�;g�b\��yFVZgc����ӻm >��]�<Rr�6^izH��:���k���Z����P<��f�I&.$Ę�O+���r8���C)vE �����H=��-^���f��OE	I��݄Lĳ'p��Q�Ќ���?4�5�
�I$í�|����X6ɤ"[l�Οc9�U��� �XG�"Iu.�ėTg�&"��W[��e�M�H�E�������b��~*7�	�8u���^9��X k>���R���g�/���1�S�o}C�$Ɉ���Vm_D���v����e�3�"ߵ�?���U�;�&�Bp�.։����4[0xM�O R���m��/;.�|o��N��HYR8���]��m���q8Ԩ��S��%LWnDZ��.�/5X�Kh��ڄ
VIg��b��{wk}י�-Em����ð!
��CHz�U� �hy���@��߰T�3�������u[Q*)���*���	B�K�|��{��[L����)��%����ǋL��β�ږ3�r,�φ[�q�@%�8����6�s�6?l%H5lo�܋�ӎ����� ��
�Qa&��X�Φ�Z�It�����$��h�F߳nwb{4�K��L�����Ǵ3|z����1эR��JoU7���#�D+2���F�M�����3��M�$g����M�z����~Z"}	P��c��bk�Yj���ebt�t:F��X����T]|��78�H�ݘ�����c�dS�;��ly'J^�J'e�L�!�&�vz���;oj"}Qv�(*�h�z�^��bb��֚b�����0�Ӵ�d�B���p��r�(�c춈�f-�!�Bô���%���w��7�P��y��5�U�ʸ�B�8Ǥs08���0�J��� �^��^p;'��[�%�و���Y��C"�1'(���۹c���I��Ȓrmh�;��H�Y�[kCAH�q$*��f0;�Q�&wE{�X
����g����W#�����]�w\}U�I����Jg��$��&��5���2
�����<���\�'�`M�Zb�| Wۜ�L}���
)�$�db|?0�dd�J�7s��f�S���M�A�����+�Q�H��E�&m�1�U�^���� mP]��f['�X���<F%ZOZYP\U�B=�SI����k��a`�.����(�z��͏�����*zEر��
���u��T��C�����T���̹�ڀ���9S�Q��������K�:k��8fN6�O �����;�r�w�U�L�Ӝ����^اBW�J�p9��>:����r���봁��G�ʗ!�=�@��r�GnA��[\H�AL��R���ת��AC(ُ�]�=���[����� �7!R��o	���+=l���dh���:��p��(+f�³HtŲ�:���#l���c�rBNk�̺���E� ��MI!A��|�V��;���AG��j`��o��͚�eY�L�k�N�K��/��7D�+��kѴJ��3�b�v�����S�`�YC~3`������%��.oi[�q�} �ƾ�֔�LG�׳���g1iW-�g�a���vu�
-UQ-ڿ���Ф/�%W)I��KC���g���Y�C���P���U�=����YC�F.�
���1��_�����g���t���g\Z���*=
zP��9zB��| )�����������8���>��uNi�!��'�,��8���5LN����[ص�X�C��XCb}�c#�9 �,ЁVv�;���G�z��S����#�@� �_j,h�7�SI���V��Z=�!���3ߎl�Iᅍ,S�@�{e$��($x@�M�[=���"3jF�&���FZ�2�NZ�3R}����x�R NWSӨ6�y� r!0�!L�2�}�����>O�V��p/���wƶ�ݦjy�H���U;���]{���ka�IR,�PdA6��d#�	Bx�l�/^�0򹷁�:Hӈ�M��i�FI��ь<��� �-�M	_k������}R���k�z�z�^>gJ�ȧ��凌�v�Oc9� �����bȤb�m�=�e��3�+�Q�~EE���qǭ�q�]��V�؞0AX�k,��D���e�?�vG\��Q7�O����O3�.hg��!$:��t�����2���.(?��v���� ��t�1��M����d�z��\�YfM��e$��u\Z/����PSJDD�}d&��=[��Zm/�}N&@%R�v�q�G�u�ߩD��C�Z2�z��]����A4�a�*�|��h�~�^��BV:�!C������"*��� hİ<㡫���'DG�i\$�dY �nA+6�z��[��&U����/���D��J{���! 0Ð�� ���>qt�����u��rt�s�-��-�F���;�����,g���^Xo�M��ƿvIʖ0�ԏB^Y|+��l3�Ka*շ�N�킰����$�
�3�Ϊ�,� ����H�F��S��`�B�-(nW�ʱ�o��)�[5�x�}o�?B�MF�h[��gs�3����4(^��N�S���5C	\;���!v
�K�
f�+�WQ�&�
�Xoa����Kb:�j�7'���~H��&�7��Y)M/=�J�S9�H�5z9:��$�[{�K��o�H���YG��[���3��9A��<Նθ��c`	��[���־�'x��
��h�����ۖ��{���W�H;���pG�uo�1,���U��#_�ػ��f�%�8����uk�L�3��X&�'�M;��ĦL�8d˛M*:�c� !��p��b�������J���l�,d���#<�CK��=f��z'�xwƛnOt|���|	���h�Z6ď�i3�3r�JWj[R�JH)��	�n�>��*铣�K=b�^$&�g4��r�5D���Y��)a��s�q7�`
;au��ޔ�&�����G�=�se7�>i�6m� H=�!��&	�o�1�t%M"�y�"T&1XU�^�;yd0��ٓ�vC��	u0�����m�䂳_��[^^H1������)q����M� ��P�8'%1���6��+�F�֟.p����2ќk�1��ó���U��1����Y�u��O�ț�9�.c�e)z:�O�~s��M?��1��F�Q�����I���Vq3�?����aq �;����t�ӧ�]F��y ���xA}��FIH���#��:\v�Vhi�]P������'�ޗø��Q'� &� �PeSI�C��=>�<��/�+�vD��6Y�Cs )��|�Ȉ+�g�2��CXe�"��~U�n���M�@	��M����Μ�1Ra�SJ��}�?:��%1FU�En/x�+w�{YV>�yD�Y
Z]��B��R0J��$y%9��"q�z|��4�C�a�I���6(���Q��h � GO5�n?�f�4�RQ�p�� ���̚=�pP;��ei	�T���2ލ7����ry���9� ������H��-J\sU>5�E�sm�5����~ܭֹ�U�[�&��פg�Ij$�����H~��ƽE��롎
l�7[�S1K��x��m�|;(t0�<�����{�Y��"EG(�Q���UV���X��m�'-P��(�����;�a�N'�:M��H��wtk9T����"	� �^!����MlM�ƛwYƗ��Ro�N���A�� </��0����s%o�}����4�#{��2T���h�$��Ʊ�_#n���85a�����D6B��)��,~%�4�ɱ�a
z?��(䩑G��~\��s���͑�.�2�м� �%v48��~�uO��`Au̮G^x�r�?Z��v���g�H���@����ࡘ�L���Z��{�0Zj��p�?�>�G#FD��P:u��*���[]N�k�
vآ��oE�u�MO�T�9^a�7����+Ii�� ��Lc��C���vqk���n��AhZ:=����������Z6u\���4u%B����&H�bl�y�
�,/��*uТ�ژ����T8!�?����<��D�<�����]ᢢ���!�'�(�Pk�C߶E���_��E������_⺲��3�N�L��R�	v�-��i��Q�R$������o,[V���Du ;�z8��Ws�l���]K]^����bM=%�3f�Di����a�� �L�\<��*	��@-�_������r��7�JQ����N@ܡ	
2ӺM!Df���>%%�����@9���/��5�j�oCs9���vay1�ϴ����q�����C륿�fc�����E�`�uo�|
eA�i-��;o��U�9=:Fd��P-1ZH{�8A�A�y?�E6J�,�����v3%x_~]��O�
����H�ac����z�Ӷ#^!��3�㾲䲲FPYȨR'�˷�3�N��X�K�Cڴ�21�M#���xY9���T ܟ��b��e' �r3Ȧ�ȸ�Fj<jB]
wzyq/����w��aa�L��`Ǟ����3��4�$S~M����vG2�_E&��9ID ��W3�y�ՄY[�~��QL�#��9Ƹ��R���N+�+�+�Em82�p�T;�?���Vy� ˬ�ra �h��m}���ڷ��;�=eRmGX�~��n_Ś��$<����ET���ޠ"G�G̝�S��8/<4e���!OBEޛ��z�_o !�Rz������d�W%��x��WE	>g�$�l=x�۠�C�(�Z�|�p���H�S$Y�n�\lg^�ī�2��x�eQ������Lf����2}��W�祭c��bR}
]���#���p��d��lj������p�(;A��=(�d��R�t���`�G�.A��0&s��JC��Z0��HBЎ�K��v�_��A���PE6 �i�"�a����@��Yu;���6�zE>�`�3�<��o'�Npaz����T~ů�<N�?w�����\C�ܧ=�h���74+Nl��VI�U�	��)(�I2w0k5]��̾Ԙzt,[� (V����}�Hz'�Ĥ%�.n
�_�Ӵ,Z�b���g>Q>iH]�p�ZV�R��숹�d�X(b�I8̔hpi�9�0dR��5��x�ԣ�t�����J`��Ϯ�c����lR��=}aC�ч��m>���6��7r��<��|Ti!�?��F��G��������d��>⶗S�� �hp��Ќ�m��-���\3������6�r��{'kIj�%8�V�4����N1�&���2�I?���ŕ�/�;I�Q&`-�'�!����\����dC���C,�(����^ʃ���!��y�%Uڧ�h^��U��}}$"���X�O���A�̡�Wl�ǖ��K*py�[et�`���J�M��ݢ�Xw�LiV�Y
~m���w�8�J�,q���2�����о�]�l����ޯ�(���nP�Vl0pI�K��joU������i����<�/��❏c�3�PS�9h���)X7@����nl�3���Vؗ����/'���_��N,�Ҏm��C0��Θ��9�j\:2�e�՜��b�4����͹7��O�ÓW��s,_���wU�Deշŏ��
č;����M�����;X�����e\u�C�Z k.G�Q�\�z�-C����{�1�Hu�̀F���^�p(����`kJ����$�/,��K��YF���
=� 1�V7�}fw��>���FL��ə%�l��Bo'��9�N��%=��,0�؏!a�2:��fN<"Y�/WԧqŶ�Il}�61���q��gj�J��1/ɷ$��Ӷ̏ �'3�!I!��P�eo��ȋ���J��M�u��dd|��D[��]��r�F�|2��u��,Z�zw��]$!iSX�
3�+؏J�'m@� �W�}�>6(��TqR(�d5�TL����`��osVtZ�|_+A�M�suOY7Q��1OP��g7te��Y��='c��o�ڊ]5,$��9`�����V�=X׆�<� f�.&����S����zy�@K�>{��G�)�PŲt�sB��Y�tY�~����O,���Q��?:z��[O$�!�M�!���y�H�u�����($���UpT(�+%r��;dj�3���ӪǽZ84�L?ᡗӕFmP����3�qAo�B`����,T��d���蠇m*Z�k�8��
�� ,%ނ4��Ѵ�)��l�8O����j�1+��t��+,��/%E�+���s�d� o K�v��cGt&�	!F�(v�&b��2HCj��kuu�<i'�\{ݎ�=ud啑g;G}�Ns�f��}@�cI��_��MM:�d+M�J�%�(���5��;w�6��(�XϲHP\�����C^_QcB݀���py@��!�͜��=�*xS4���spN���r'��r�C�TO�%j_��?EiN����R�0;(2�GY��:xazNX�/,n�R˦��;�R�A$�G���8�L���{�(�}��iMd��i������.�����w�`\�L����"��I0�\��29�y���+#���)t[�#�Q�u#�ߒU~A��Hk�Gǧ���\�{\Zw��q#=j&/ruU��s��Qi�D�au8]�"���4%R�_�a�특AW{2�;a�F��WD�K��`}��;��V�F*vW�K��O��?"�b$c��
[
������žQ�^�^U�i�Ѫ����?�ֻ�Ӧ�n�𐎈�36���;{ƕ�E%c�+�M��i�����Q0õFx�� ���u���|��-b�M�L`H9c(ϗ1[$齉.I�˽|��v�l�:�spW�K���V+=.�=|��ot���h��!1aZ��[h�-2WDVn���8�e�2�g��nF:t�i72��Uq�m"�iӕ�7�F��]�s��
�uK�[�\"˾���h��c�TN��6B����oȷX�$�=�R����_x"9N�P&	� ��reuc���\�M&m��k�"Zwj���q92���#��/���L�>6�H���,�v2R��͡1�73� ���a�L^K'�1��//�Q򘬦�\
�I3�b�Ç<��&�c����  Y�$j�hXd����ʠ
���.�H��G~��b7Dk���V�}��e��w��[Jc6��X�Z(LF����A�c�ey��m	4j��sȮA�-ޕ)��i�?�[�H@bK>�]s�C�2`ɶ���X������3:�����T	���5��>zO��.�.�y �}y�ed��{�����V|��{�,��=���|c|�4�P����wl�ʔ�l�FR{��N��#��hJ���-�?���K^����%��b�e �j��������5���c�����t:��fz���p����̮4�ʜ�n�`����G��1��J�� �D����,}����͋:|��ڧ�3(�>�93J���0�9������n�McK])�/@���O/�N�� ǧk�zK&gA�_���-E���l� y��;�d�W�i����GK��#�4���&���`�Rt���x>^�f�]��������sDJ��sS��P����A������o��I%}eVx���L��,{ ����Z����\���8t��fB�y���@$�W;��~NS�)��(�_�%"ܕ�Q}��^��f	,a�HШ����皢��&~���`Fv-S���~.�[#h�"�G	�	������r>�	
�5��K�ո��1r��������|G�qp����+���@�Z%�K��p��~ͼ+ʑ n�~�G���'�IAqKO�p�p����=����
J�Ռ�9lQ��j��db��b�e�؟�~I� ,)��a�4�����Ȥ�����ݏ?�����6p/����U0S�l����6�t�t6��Yu]�B��#�]�u���UQ"�ß�OM�$"r����w�'�c�Ыe��Aڨh������O�n��/����@�>�6��'O;@�E��,���ۀ �T��BF4>3�uؗҵ�'ne�dgFcȁR��9�Ӆ��R����Ĥ�H�!�:���Ke c3K(حz@���i��6�k�M{�ȃ���X>bU]y�19S�}��!�+�Y��^fu�ih��Ɯ�����{9^�2�
�
��E\c��:MX#����;����(��+\��?��>IH%@@Ĕ�k���1����q��� W��}*��z=C!,Ǥ�G�#�_�HĠb�2��oq��M]ĭ����\��"�Ą����ko'J5+�\���e��߲$�}(��
b�	owN�gg��-�V��˳��yi]��+�2!�͋���XN����0��eT V\�'��u)���O�"e����פ	�l�48�i��I�W�(�}3�h��~X⨴�F�0��v�F����8���L|��WT�M~�o��T��{d��td�|@��iMv?D5p�$�M�~�j�����+	��I��eP��P��0]M�����+�����<t�ß?�:1n*�Þ��P6P��d?�Mp28�+�Ot�)�~W����L�>�����	u��5�1oC����v����+d��,�N�tc����9;q�U|8L�&�t�{�M~o
��Ab�j�vx����U����r���R�cZ�L:�uq�' d\���1CRu
;��/k�[2Ҝ�A�=�������_SYW#���_���?������<KPy����M��m-5hAs7����J��k����q���
��h� T�#�v�R�b'��Љ
��p�m`g����T3����Rzt�ho{`Kkd)���zjJ�m%��H�7�q~��zy��@��vPǦ<J�1?��ހg���dٞ��_�q������K�W~ЕDP���^T�)3�Sd7��tY�rU;����$�>I q.>S�����|8h�	�?�d
fox��RytUnB��I\����ww�NQ�`̈;�Dni�{#��~=��b�"�p�/��$Zp��{t89"]�7���V�?)���y0�%%�+f�iO�a�����k\�1��ȁ$z(6!~I<؅�,B�v����[�ERW�
\��������:{��C��p�F2	ER���5'u:��$���Tiʩ��w��L�{^a��3l6Ό/�ڇH��.�A�T�m٠o8����r̹�26QCF��䴉ފ/��H�t�ΘO�o*��{$��͓<�y�6Bw�q��C���	A�鈘bmxa31qȇl�yS��tQ�w>s��c>3!�;�Q�pY��
2�%�
�̰�/�f��#@kI��8�
{ܓq���&h�%e�'� �0�4�s���'�'���X������]����_C��=-���CG�XY�f\��[N	v")���%z��%�&���9���3a��R
���Qm[͈�U?�/�<�y����V��v��5Q��{�	<>S���ɉy�Fz)Լ�G�x���#q2�@�R|���-O`[APL(dd6����Hab ����9��4R[��e�&A�]R
9�K"�6oG?��� 
E��^q��pL���V�k7��q�f���<]���jL��DgK��ӧJ7�a��p|P2;�`$��L�)�cM]<��uI�,��Xq���hz�>�!/<����A�8��m���n&C����~1��z�oA9J����7�s<}鸱�^$��)Cr$.ϸ��W���j���X֐�dQ���}Y�7��Cr�����o�"�W�<�������
м���ۆJ�jyW/w�l�T��o�g� L��yEȮOy��Ɣ�G�RBҟ������'8
c?���+۝f���C�bˊE��
������h���k��A/?�[R(�� /�Q��I�Βk�NӤ���*#�|i?>�����&qp�8�C����Px�f�~��\~X�O�K��0��ſ��8Zz6�Pa�<o�w�A�:� ~���_,IWZ�оD=��7�.٫���X�[�+���(C?,��ò� ���'���&W��5;����q�1D:R��A�}���N}ݖ_8�I�SqI��V����{d�F����ge��Q��ˌ�W=qc���q�L�-��V�7�4;��8U���{9�q2@�N6�ײ+@���Q0���#hò.����K��A�K�\�����C,l��Ѳ�_
2��l+�Cm�0����f�]��'JB�O�� ���L�p�F�M�<�����d�R�:�6`0Tr�ĝ�4x_f�R�&I��E)���C���h��*/�R���T&����Y�	��Ǝ��hQ�����XP�[�T��'���=��`o9�=�S�@ԆNa 3$�W�z&�j7��	hL�|EU{�1�S�a���Z�,��hp�S��ju��g���d��1Ź>��jy��q�3������2����P;A��@ϰ����>�gk�p��|�c���*<Q49� ��ص^�֧���t؝��j"��^8юP������y�9�v�R�A{W6���g,��b�O�=�-�ֵ��>4�6@��y|��P1�(��g�
c�И������!�}�I�@I���(��>�����ʃ߁���˾����m.��Mf�S�iݑ��`a*;�	�|Z��&f�럖ǨOx���,�ʽ(t{�x�5oO���BYU蔺<^4�2�Gh�
�6�M�[$l�X�5Мā���(! �[ﲡ&5���!���aWm�?Rΐ����}�������k�!��������p�M��,s~ r���Yɱ_&��1�L� ��?�s�]6N�U.�]�T�2��g\��8q)#)�\�C"���
}|2����7��!-�1
�#o�F(�'� ˂,aߢ!l�߯$��ƶ$�%k�5�]� a�:�g�N.)^Y|�$ �%�8<�lE���I�s����^ć2�>�W���|��׭�n�)�LH8��P(��;&���3Y�����<M�X����ãs_� jV��� �u�& �A6�\��HQ�,O|S6\ϒ�20�1*����Y,K��2���`G#c���|�o���N�:/���Ӊ�{��x�����a|����׺��r^�k���ع�8p�M�a姦��lL$���!=���Z�6^z�­������d��3��Ac���տ|��*���&�!ǃlb4�/3s>x�j�Z��7����QÅ.�ԍ@dI�0�x"v_��<�]�[�&|v�w{&Ț�Vql|��Y@I��`���l����K�c�O�z'sQ�cH3:f�L����F*�S��� R�~N89�@��ľ+m��xm��	;�e��b5',���ۤ�G[�5���~3��U���j���R�x��d��� t"��qsHM]��?�_��"���sj�Glz#�EQ�/���>����OH�%[���!X���$�fyӟfP�"�~T
���B������_�P��S�/#�X�6�Z�ZH�aF�����r�\}�n/k�bY�Pq����'�bh�v֯园we�q?���:����'�0D���k�t�Ӝ7�aO�V�E�>j�<���.���5�_��y���K)�v�����䋤k��~��_g�o�ʖSOv����P��
���.�3w��7mcVMv�|-Q	���t�ha~8B�������)��|-	V���>Āϕ�:l���8\3��?h�s��Zt�m�3�ƺ[�7S��AF!��7!
�� �.���KU%Vʄ�� �2
*�q�H�\"\��J�j@��i{)]i�վo֕������P���Z7���T
���F��?��|���hD�:פ�_��B�쨄i��4�o�+>�1�3ĉ�,"�lF�$C�b�ȶ.�X��n��	���)��*�G-۾EM:0�(n�@�T���]�\�~���u���@�j���mMi��G|�N��&.yW���ۄ�N�S����R��n�	C|!�8?�l2���p5�
z;�eRU���hZ;�FU���W9A����d~P1�\Kݰ�̅~~�>�Տ���$|[`�n	s��|wq�
#��Ie�>��`n�D�������>�Ɵ�j��n���z7V�g߻��<ֵ'� o|���L`[5��Z�Nu�����E��J��^��������ݚPz�8���¡gs��ut�&�Z����QC�^q`8C	!��x���La�Mf�:K��0 ��;q�75^4g���DI�b�?��s�8j�$�(�d5`�P��۪a ���F5t.{��7n1H�³�]���v���['&��<'� C�K���c�s�M�\�^i�y1�0->�"�8�x>]�T�&� P4`Y����*`��3���c��}�#�-��cc���&0���/�"���˹��:%�u�Pd��hYb�>��@)�na��,�=ѷ�-IH���\�܈ͦy*Z*�xw�:�91�n�v>Q��M��t��O���S/t{Y����2ЄMl0x��[�n����)Q"����k�,t�<�R7�7T��|2�fv&~�O���~��@������|�߾�7�62���$����
E�M�c�G�V(q�\��}fɓ�D�v���A�֓�o�_iF�G�`�]Ro������jL���3�4�rubA}�׼�7���O��)mi.�_����k�����.�nW[��e���L�S�����U.��JŹ��Ý�x���!Ԃ�ۭ��?Q ��"����t�7uԈ�g?#BY�%�
TA �^d���;�������yŮW�J(�;.a��\���w�\?#�����#�1Q�J�F�����̭���@�"�^;(�l��X��f
ZV���~�XԎ i#Uf�܏K��p=��x���� ����V��L�2{�k���Ȁå;����O�:�5����K`"m��V�3�w�ܻPH�.	+z�Td��OC�ܛ~��%W�zE�����zM�{���R����/��C�uՄ��<Tk�JWF�`G{^��Śc�5C.��>�vm���e�y�H�k�ɚ&� Q`|FZ�3ڄJ1O��}�X��tl}S����XB���q���1���]^@ޏ[C<0��pVQ1�[<0?�OkA�8��)�ݛ���(�:�[Y�+w�/ �� q��#M�R޲��kj�������3@�[-�w��A��j�zVlG��_M�Hqay�����ՂwC�b��L��{���he~�����B�<?�1u?xzU�Ϋ�-�lGƗ��#�����kk��孻_�@Vk��`2��g0���Ԁ��ɮ*�bQ��2�W� ������DiA}�n'Cf��|�f�=8ȯ��<��6X.���j�ψ�D�`^�CZ�4���pMC�
(��&�/���oύ_���vp��I�-��7�%W����n��&p4w4T=pL~w���Sy��=�9Gj�����A�#�M��;^�2��:�{�}���ͅ�=��{�)�t�3��EX��sB=J�bȄ����-*Ŧ�"�Ք�wLm)C��÷�������T~uB<V�Mr�L
��u~��-"�=zS|�!�W-�,��ʌ�h�F	_[��+�.������t�W����'��op�*��4���v�������T1Ҋ3����߰{d��G	,y�r~�'�!{����{����U>��]��ݸ卲���Z���2�\!���rP,� j4kd�q"��'A�R"~�������7v[�A>�S��^
}s����j)�b���g7���@t�ӣC�6�S��&g��7�P��m�ՙO�]��Y��|�b([��ua���>�l��Ҷ:�k�q]�@��#�o X��S/e|��Ў���e��-���[2&�T�&[@դ'�	��e�%���V8 ��(.GV���2���$�o�}�p+�O��E_��{�d��'����?�@钔a��!�,�.k�mvZ��O������_.��M֚cE��I�v��ױ��v�c0qmKSS�Q:M8�6��њ��<�P^<�L��1�;q�.��j��F�+5����ٙޚnXL_?�o�$a�����?"�����~E
��,��l�0&��䇡6������J����Q��Ӽޚ��D�L�� �	<2�V�ë��X_+��]��b��>�JP|�g�ep%#�zx�:�D�{b��B<��Pc����T ���u;an���7,�f�e��e��H��=�/�6���&��QA��h!�=���f�;))
t/�g(ܢ2@e��c��7Ppv����o*T�on�.�^2L[J�_�&p2��8�n�#4�0�{�O��Ɠ������"GÞ{q#�';Q���AjQ2+�A��Y�ĩgTE13���ba��Gť�]����6 Y={ÍX]v}I"����s��;�}��2:���%�a�XS)W�QZ�^ }U��tPcU�Fu�[:����)ZzPD�m�0���4~X3�	n4�)� V���l�(��H˻�<�"_��u��9�U��?�����|GӶ!9	:������Ř�Vm��"F9:�?Yc����4�!�4��"n6�	���?L%|ѿ!�"6��C��°��?����z�3��W�p��I��~r|�S��M�@�Go�p���j1�|�/i3�\iH�!��O�ߝ�Y:Y�@��ɖ�|���!��P�}�H#��;*AH���*}��'�#�Gmٙ>����<����g��X���X�I�o:,�Ng����Uhe�y��|�����ػ��L&��B�T�{�X}?~-6bkEZI�;�T2�Pb�&��0�L��C�ߓ��H+fh8 2���´V�ѭ?z���r�Q���a���_]5�"�j��u+��K�8�:�;k���D67�=��̵ъ�च�I1Y���ɪr�g�F��OP��
�8���*nUnt������.���ܿ�x�b���<dɦ'z�u�5C��6�a+�+�E��<3uUZM�X�}X�����}�U�7(:|,���j�Կ����0�\�t\�ٚ���f�;-��!^�o��K�+���o��O��#�,a���� }&e�i�p�9p�W�LՊOJ��!������*�J�9�*�c�vf,m$a)h����	#P�HID�헎�H�N_F�����e��$z8Ӣz�8uAUBK^RC��H�ڍ`˄_��h�|`~����y����axW�;X��h�~������!R���Ӂ�c��oL�*ޢ ���"]I!ƎCI� (�E���� ��.�y��N-���^D�'͸o��ۭ����a9i��N��>��ܢ����b�0.�p2��T>͗���vuhjƨ���{o���2k�`��'�"�?--C��)��a3�2����t��i�0����{�e���m���i�7dLk�iV7`B����Hd*��.Tt7������
V���٠X�m���;�K��K���_E{��9�X�ǖ��=W�]�K!�`���65#�����Zgx��3�VPV�}7�1�� }����̅'6�+�|m�BE���x��{�/���%H�9IC�i*zB�~�u��Z�G{cW��U��IoB�k30 ~VðM��_�,�����%��X�F�:���NX�l���|f�0u<�<Ė�7b.[poBg�p�,ٺ�)㕴��-�,����.�x�*]�����`QqTw3��j��� �`QO�WL>�J`�u5p�NUQ�9��1��	ݻ�+_E���
D��1��TrS���5E��D+R�IrO�!��_���$�����ׄ��Z�>�Q��#�����_�&<e���lXX�d ���uw�ߝ�|$������B��Q���5��+R&��ˬ�bԡ�9��B0k:}W���Ƌ�F5���ޝ�a,�T^|�ќO���@��Z� ��:�[�#���Z�O#Z��AѢ@�)`���j�T�O���nC�p���6WvVPy}3�j�/�@ �a��SҪ�mL������M��>"�'�
Snr�����%!CԲ��%�F�8����$�����eP9W>$�����`��l���@�Z�(�����f��;����!�p�^y��gN����Vtrr,y�$ۢ��KoR� ��"!��s��qCN�c����RZ�9�b�g2�_�KYc�C��ZD�������@�Sf�����͐�=է</��2q���)J��2���d�HJ] �?6\W����JK#�t|�����,U�]?�t
R��IfsU��!�'��n�gt�-���T�|�P_K�{��b��h�{�Q�GR�am��}�U�w4���RP��~0k-��l}��k�H*O�����#��$�����9Q��H���>�?^9W�$B�0)��5�]H�ꇟW��a�E�լ��� �,G�0Q��}�����:)��M,P�� ��4���4�ތ���-�|�V���@�w��ZB�k�������e2�_���!����R�@3�ɉ�O/��qċ�� u�n�I0��{H� 1�j�cO���Ku����S���T��ҥ.g��,���&3>�>󅿵 ����r��"�]UѢ!�2Y��DV�na ^�⊊���O�p�7�Q�=������������v �E��M*ri��jb�q���w'�����N�k5:�w�};_��+�^�̌<"��j�(���ͨ���Q�TM� �<ě�~���"�Vզ�X Ă졏fY΢���K�T��S��d�>��hi�V��X:�;3A��m�I���y�@-�;0M����Y�vۑ�O�N��ow ���}Hy�1�ޘ���scM�`�c�E1n�e5���Q�F������꾵*��P|3��#w�	'0��G`a8��= _�8.�5�5��M�S�r�4(�k� �k�,p�DTr8K����<��ՌV>$Z2<^�5�F��Aa4.�u��s���ˠ	��ƫ���"�`���GzU�������*�y�o�/s����aj�U��8_d$߶v�[�����6�/��a��^�r|�X|� ���^E�t�Lm�Y�l���:<�tHΞ���Q���,/S&��>f�Y����	���7�x��V��Yj���gt��b{c՟����.��]�r��Z�����^�-����%>�U���q�dI�7Z�}͇Fȷ+�r���U7���h׷_C��!��7�-Uu�X���[��~-I��(^�XgO�(~��&g��Rn�VS0�J�"K���q���ZX��æ�I`�ˀZ�ETS�Y�^��W&y�4����9��'[�,���Ȥ���T�Y��!$/V�;jK�x繵G~o� �@
��P7)q���E":-�Ƀm�,f�����|��$g"4s��$i����~>R08��bΊCR�R��u�b�d�B�oYIQ�[T�cpb@�a�!����KEc���zؖ7DN;���Q2��_��R8�\acBuk\.�_�a[3ϋ��ns
)+����Yh[���۷V���~���)�I�W�ڢ�{r���g�l�jc�Ԕ�r��X��>����b��MH-Ń���sU�Hw��p�?�"��*+a)�+��MX��h��Iq#y@� �� �Ð�V�IWc�<kg������Q���-r��L�~�ȹ\W��Q��F�G�Y�s,��e���N��
0�E��3�}���������S��\R�ӏ������N�+(gc<!�Z�
8��Y[�VM���z�l?�)���&��Bb�%�>a����	jJ��߼��q�t�n��(�O�g+y�:Y� �^5�q(�@�G���S?��p���?���4�=�_OV��|�)[&�����1�6��~(�ND���9��%zF�FH�l�?���`
�����I1��˝>6���߂��Y�I�:��´3��'�0��ݳ$��8n�yBy���q��|�@�_V�M�����$��t�x~!{6��;{,�;x$�b�4�P/gv2���X���\_|G�^��lB�X���$�!�����~4sCPb�A��Y�$+�T2�:�cԅ��Z���N]�h1�����ݥ�3.�S�;GI�����I����#M�,QW�+�%�g�7���*�2�0+�E���{4jw�nz�~̂��o",��7h�u!����Oq��q��^g3yJd��k�>[n�>uX�W���Δ�
�>��_'Ѱi�G�k�ڼdR���AJ-�B�3�7ʩO�Z[�����/{�F����<���u�mW7�7z���1�F�*;�3�qA4�d�\���u-��q�w���h|&����H��ޢ�KyKH����8��M�#��݇,��f~�|x�'��E
r8ԍ���OϣP�z���֭��>A.f9ο5=�1ۈZ
�wR��PՖ���m0Dy&��){x�,�P�� �ِb�9苒*:��OZ=�#�-t*1�CkJR.� ��N����&fٸ�A�Q��>ړ�g	n�I�ZQmd�D�&��[���WH���9�ɨd����X��,�2\���	�фV��c(>�X���Wی|�����L����U?�����:ɬT����$�f�������)ц���c��=���[�� ��vE��?����D�]������c��<��E7�yOp�]}]tG�3'�)H�\��;���"�L�--�Z���?�xc���{��`�fP�t�$���QQ�7�A�� rޚ֏���:�X1� j;V;c(E"�=*�~1��ٕu�ܸ��Y8��:kP�0c37�������J�弾
�P�w��|4 Ug~[�z�)?u�+O�x�NΡׯ�U�8W�����o�'����0�?�P��9U#��a$@��.��Ǫ�A���PJ:n�*u9a�+r@�F<�p�4k�>�wa��58%��������\
Y�cpC�̟U�ne��T��׶v)T��$�ʁS��X܌w�`�uۃ�^� Y�|/���	��ިŽ�U�oX&�q�<T��<���� �G��b/`�.�/����h&R+���1d�-_�R�H""QԨ������q�\F��Z	�?+���� <v�®Q_�Ӿ6���P�֎�B����B�tt����" \/P��aHȪ����Q��e�t�	W��#�Ҵ��|�/���'̚5:�Fg�`����Q̸IM�]���[D9�f�v���Tn�|��ڛ�]0*�O+!�Y^�_�,����6�_�OAJ��e���B'Wb�!�=%(��Sw��5(aAȘA�7�o����p��%M�U�*=~�ۻ��R��:]%0�V �;'X �T��&���������o@�����N�HX*�Z
��y �1ח�¸�*7t���cP�q�ԍ��U��c�����v
YR���	[��ɄX�J�+9C�ӄԿI�����?��NW,|W%��W-v+\��5��U0׍��g>_�����C�`����C{��ާ����� nd��/�el۞z$Ar�Wi�S��uX��2aX��ɖ]S�6��	~r�/��ˬ��S���Ez|󎎄���d�+��=�p�%H0�]���qBs}<U�n+�[�Lپ�k����}x-,|+}�0@�W)�1���h���r��t�ƥ�b<��ĸ����ei9(̣�{q&A��fo�4N�(Y�u��M��F8̜d��D���+��r`:�[��1Bu�[�G}�x�����ɥ�?�s,�lph
w/�'7\��r���N��
�!DރW�������!�&����Nr��F~�Bo�������ja-��:8�	�Vyf"%������� Y"-��ƂR��%�.�����ypC�>M�v>���th�#d��A�2�(��`,��S��wNr��8=FP��[�@��%Y3����T%��������ܩ�eKeKj�3=L�0G�z�WϬA <z��5� iF�`R�(]�tDD���!���:k.B�&{�ձR�#?QU�7�"ǂ=Dw�v��c~Eb\0E\C�,.$���f�_�=�����Ge"Ƚ0��:��zW)Jk�7u�c�*���&$���E���KL�Y8�ņ ;��ˆ���M��V
�\J���e) ���I8׫�����8���0?��E�_Kh�r,�0g���k�׫cs��@) �#���S���h,׀���N�c���u�9 �^�4��d�{�'�9^X-��7��
��v䴲xYC�Q	3X��΀=C�U3 cm�_��}\1#<ؖz�4C������碻q��5�Z5������ ��	,O��;ŒD#�G���tA�Vץ�]G�(�va�Z�`֮{���bm�,�hu���n�g3����u�7��+{�J�6:	j���77>$�|��n�<$�4S��[�����s�y�IB�a�x������]�a�t�BL���T>.�*�	�-���j���	Eou>7�8� �(~�W/Q}u(�K.\=R<���G�n����s��Ğ>��ũ^�N��b*�T�a�z�F��&�28#N/>�㉐٫��tdm�l�G�2O�vm@��uA����,������X���s6xV%�6frS��D�<s���c_��d�a?���Zm4a�v1�BCG�������Z'����Ҏh2�|���m��=r�N��I7v/vG�K���<?���iFg�~���8�G��ZY��_�o�i)�C%��~U��r�׫��%X�Z.�#V��ښ��?��H�8�v��+�g�6 ����|��� �4j�~I����J�8٫-����Nx�D�^�~�'��^O6��=�F� ވ\����r�����b�W�;�s��]Sq����/&�)������."�_�F"wu2g��_�$L&��-#��m�A�D}��K�yc�h��BU̓yO���n����B�"��*�*������H>�-'$;&4�mի�"T��al��Rﻘ���κ}�^d0�B�C�(ķZ��&H�C:P?#�9}����'I&ɘ�������
d#z7��<������e5NX�j��"����ĵ�Fy�܃�=�gN�)}�$�tVo�l���(�]\-GY?��*7���i��J��U`-�&�����I����](d�T 4έ^R�������7Y_��;��$K`a��!�3n]��5��������wR����y�\�~��^�{���v�G��	�ˡ�C�_���=7��|=u8M�|N�1c���E�l�v��|U�����hy�� �'CQy"�Gc��s?�j�6�_:,�/�eo~u�q�b?�V�D}���96����U�����{��4�Ymo'����̝3�s��μ�%�UPN+��%�j!�/%���#��T��_��m�]�Y+/d�R��js����k��"����JgT�%����~�Z��c��ы�3Ѱ_��E^��
��L@"Y4C^�}�������8�/���Z�i��Y¬2'V��!�GF*� �`�p �D�̝ҥ�5{����)W�	˚����-���h�͓�c
�#={�|�z���A��K&��?���X����	�����r}ܲ%$ק,�?�l�#��H�5,�V���0���_�%�6݈�������w��M�K��E�#�tk��� ��3��}�;E�P��(>��	c	g�$�-,8���5�� 0,]�e�%���G�Wa{��Sz������Vf�U�[1?�r���85#��	�m�Ve/�+b 9O��^yfV�t0���	��sƻ5/�����>w�P���~��M�&�$ҋ���gro���{�	g�t[ꗯ���؏�����2����G�Zr4<����g�Ψ�������T	"��ɳr�Ow�ԝ�22|����ke�?C-��y����2Æ{��y/��ꋽn_ᆩ�(�*fIϔa��~ϲ���)b����0Z�U$z����B�D�#`��jgI���`�Oīw8C�?�����93DM}��6���%���0�{� :��<;B��ɦ���x{�>yE�����C�V���c]�>ė���K��o��A���G<W�8I�ҟ�@x�7	���S@�����R!����\������ �G�l��9!OU�0�iŵ������G��G=��@���(����k$v����	��C��^�k�������q�
�P��&Zk(�r��x�4t�"�`{r���2n�������_Yΐ��������
e_�e�J��O	��<�C�s��ю����΋~YK֟�ߊ���VO���Hj��}�c��f4����Z8r�^��c_S ��M�i�*_��mGM#�h:3�m��:�h�}�J���s�E
�q`�e�K��]��Sо��	zO�J�R�U���>��iS!��]K�Zʯb�?�v��T�f�)_��Z#�	J�<1跦6�ef������� �	_uk���m�5����fX����G�v ��7~+�[���S��ˎ���w�QR�'��0���Wf�ǳOs��c3��@�ct�޺v�&LE����ޯg+&{R¾�.ŉ�t��6�B6��������M�z�f'�ϩ�7�(�g��òa��%ƕ���®.0y��X	:������vzD��g��aF>�	9�9;�&�:�e��cx���^��$�r�E�J��-S�����H؍��_�O�9�Cr"~p�43��ᑁ]���N��_�0�3�;J���9�� s����Η>��7�t�N��GU���-��+��/f�$�R��¿��j�F�dB����#�" J҂�+�e��S��{'�Jhf���Rr�i�}�׷���Լ2���ⵋ�5�A�
^ح4��ΏX��i	bg�&fU8) ��-@������s�
a��>�*��b��!��Ec��QT�Ά�S��F�r��sJ��8<#Tz�	Z�ޗ��G�aQ����B!�/�MwPݕ�f#�<q��v����4>��g��SF^�zY*52T�b��كe]t��RP#:h����p d�!���ݫLs� � l�]���M����V�4���9�E^g�T!��F��ƚ�s7l��T�h@�A��;M�s�3�� F$��d�Eu���/�a�����7�B9�;C��(PO��^���!Fn��v��S��i	X-i<l�ȭ���X	h�?
3jFt6�R�$�A ����b�+4�,�B�3�E'w��-4vo>���}�_\�������0�������	�'�j0�(3a���9q{�c�Ӏ�p|��o7��d:��in���Q@M��hS���لCz𩨧�����h�av����
?�&�W�Q�+��nn[����[�[�����P9V�a�:щ���4��1&�	(�H����m97�A�W.`E�%������jȫ4�J��p��$Vd�O���3�~��&�B/���#�~\1JF��zq p�@�]ؿ/Bf9۟�M%�<:TDP|����e���w¯C�`4�T
�x�%ixG����$�tQ���h��_x�֢P@�	C;�p�y�����^���@����yp��׬�h$`��Jr�v����ED��7��� ��M�@����?Qa��gc);K󆁓Yk�p��<$ßݫd��k/��9�+��R?	1���	}N���ǋ��z���0*�kγU<�i�u��� ��S�V[����)x^�KmCr��Ք�a������Yh�\'yN�1��s9A��qr��گ�,�k�.Г]SMm� l�Z�|:=iA�2�6Qy��pz7g��)a�f�"�w�ચ�<��y=fm��ސ�O"��p��t2��S�Y|�<=I�-"8��-t��+sm�xC�e +B�ߧI`0������_��[�:������˕S�+Ξwi����OV��ih^��;��D�>�5hN���F�?D�ͩx辶� G�N�6kx�u>u��4��o7�/4"QӚ���*Ɋ2�ld�C��裭<�9f C���T����0�܇����_Άo\�dl�ٍs��\U�Lk��b�D��H�"PII��V�]$e�v�}EvԩYB�+Hѭ�8\����}��?���`�����1fQ�F||45�m�Ӫ�Y�ʝ�VD�)+2�Z�@G��P~ǚ�!wՓ"��N${��%���l��W��~0w��/G�.l��{�'Rk4����l|Ȥ. �?/^Dq�����,&������\�	�k���4����͚<+@��E�#Q�=!M&S����O\ާ��W '�2�0�Y����V�'$�6c�h�e��	��fM_���-���9�Fb��g��8�Y�8*�
bc#��A�������ـ���zv%2��x�O��x���8��T[�rv`6���<Nvp����_�����PB�����UMK���jG�������-���Vj�a/�f������!�����r�2
�[��:��#�_2c��*�������Do3O�(�K��
ȷagb�^���9��_9�4�J�n�f}W}���[`�����o��z!~�f�C0ci<�����ۡ��V	�I�z�inާr�KI�~LB���I��˓��OO0v?a�<0ЂEX���zlY4��v�W#f��aih{[և}+G���=q;���I�̲���^z���碍C+X�:.��X��-'�DȌ��_r���a��Т1���=��.h}g�)<x��^���/11^�iI���P��o2x�8��wɇd{=�D��9�q����X���8'6���%���ߢ���q�F��9+I�� ��}5�ײ����/��J�ø>�Դ:{��p��"\���=��C�$Ŗ7��\(U�!E̬�@�V!��p������^)��Fٚ,Z�����%d�@4�!�Js�e�2���� *���� �A��;��_U3��%�R�y���#Y� ��R�i����v>C�����(S8�/}!�H}A��N�/5�Y 2�V��"E�1G|``���"�Ė�*��+�G��R9��z�E���Ӌ�ق�F�g�NTo]��m����d|���ۉ|yq ���~�'Ȓ�E�ʿ��O���LL�_����)y��T�+=Y���^1%�kTy��s�i����Y���;�nA��:��x@��R���l�m��A��*|�A|�Jo'��.���{�Z�JivZfV?�^���y��R��?��%�>(R�##(%0q	oѫX�	��2m�㟴մ��a���}�0�c�(���v�;&z�X/�QM@��[��n��7^�)r�����r����">�J�p�"9��@S?B�B�Y*�>I^C�������ӭ�9W����f	ل��9s>f�Z�R�'����DZ��m
~��O�w�_���/(|�=��Dq���MXs���ޠ��ieE눖T���M���ܨoJ V��>�^����dYD�<�մӞ۔~^�)����/��G�Վ��T�2�+�[�cQ������\hJ�<H*_�~������W�t�ڦ��	M�cQ�)=7��(�_&�9ma�D�7����-ǩ(����W�|����T��~SȲ{�T�BY�����e%ֹ��?W�F�G��c�q�T��v:�������n��A��MNI�k�y9��j|7�cJ����=�{����;Y~jH/n�u�0=���^x��YG�l[����s��jTʲ���� a5����������i�F��8=���^��~]Z暝F��{~P�����C������W�I��������#>�������*�������L_ż���zhF���uz���r��Gu~ �"�.����<�q��9�F���c����`�M���V�6�{��6�Q�#_Ct����^��b}�Z��?<@?�zF�H��i޸�G��2���0wCrD�BDD�v:6��?�π
��&��f!hc'~�e�ԧ5�R���xūY~.$�9mb�����)!�ڨ�'��jL_��!#�H0�)S�����T?��^�Y7[���@� L`m�d��C_k4´,#��?6���m���|v�]*#�9��r���������w���`��Lߝ}FsH}vB��J˙��I2�7����J��z���EC1[��;�$�����C�$#��b��tI(�6]��;Z�q��"�a!
�<WA�>O��>D��X4o�DQ�V�5�G!YA���Z�FMb�|8�+$�YQ���].�=��+	*�r�ѮZ��`�=൞��x��E�#A|z�5+d�^{�Mu�Tv�Q�D�E�2
N�U=~�D���#�uV�¥U���v�/�CL��k�^u��ϲ*��LӲ���ͱ{ c��Pc&�h3�D��ɋ�t�KS`r��ڔ�w϶��.���,�v��ѡ�2���k�U��ˌa���m�G���y!x�M�?����' ���E���b_ؑ@�J����l�I�x��$r�b�ɡg�a�$g�4Aޢ�[j��`������Ԕxҡ���}Yc��[���B����On:���°�N/虰�3�>����N*cʢ2�"��2enӇ�W��e��[�0��4�p�?#uRn�����>v�
 ˑ'��M�jT��i�=�A�HQ�N	f�?���Q�e�IO���h-\�T*�,�	�:K����1���,�]��ؖaPV	���o��������2�0�aƱ0���g�)�����U���>*а� �|¡?�:W�q�$*���~a,�!n��;�}r�?�1C�'ezq�[�鉭�͚d�[(�n�5�*ژ�5bh��Pxbd�:���0g�'���\Y�8�bR��2�m�sҌ �$��uYG���C�r�)��z��'	/�?7 ��|{�b�$��v�Pp�������"$���Y	ya>&:����K���E����5��Mru�K�z�S��7H��j@�&z.z�	B�_��ip���F�ж�뒶�/Le�0&C8�۪Cc�4tI}7>��y���흔���x��v}����:�Tm^ID�O���.�J뵇9�A�È�iB�5�>��-�++�r��z��i��Q���2h}������-�z.�d��|�����_�z�-&�'����t����v;E�A:�f5)|D����<�P�B�o���ک�^5~plB�W�t�:OZ�R�w�]�<Y�s���&�����A��X�< �Fd&��q\�J&�Bk ZX��F4م����?m*�(��VIx�G曽��F�e�,�ŕl�[��k�h
���*C}�s5�z+q�N�и�@+�ޠ�x�'��@�����yK�Vޒ�q7Æ�����u�D�(V�uP��|ޡ��r�Ӿ�y�
]� �<�As��ۉ6�����]zM��+��=�3_��np�*�1��-�j#;-��:�w�y{	l���JS%��tQ�/��m%.�q#H�!e ���4<�� 1HZ�����o�7��nӬ�J�a�i��OA�g�kFfs��'���Gʴ=XҜ��&o1�V�Q�#�Y���/�b��Ĭ�ܦ|'��������}�X����uPM�}�ϰ�k'��s{�N/zV�(`q"]�P��WOt�����J�s�V��u@M�҆Af��=-����������oG��t2b�j،��I�B1[�fqf+g��?]KS�P*�ڭR� �X��-�Y�8H��6�d� ��p:H"�1���Կ�W}�r����ְ�u�f���zm{^w[6����{i�5X�]f���u
H�*b�
��W�I��2�W��-����#Sl�z���f�V�K���]G�$�.�\E)�J'V�ڦO���
�o�e�� y��-�˞�lߙ")�����.�'[�k�[�����@��fTa�Z^݃�y 4��%�~��?[�9D���o{e��Ld��YZ���Tk�(���J����e��{6��>�~�)�v�%�jz2emZ���XUK1��w��"BX�7� F���P�É������S���.瞮��G���
�.�-jƺy~�$ㆯM��fؘ�I��'�vWiauЕ��:k�D������8�ģQ���*�]x���p��c3�S �BjfT�1�G%��Y�=�Ȥ����5�J��=���a����l�9�q��g ���`*��Imz����M_#��ژvv?��V���;�Ζ�1>��^�ʉ7Y��E/�(Ù���4F,Z3\1��%e�L�N�'�����+������/@f+ÿE	��Y�䚝Q2�%?�^�w0ɪ�Kw�_�33e�.Ҵ#�H��'�y-gC��1����U@�%�5��K��{rg���tz�M��z(��u݂�r�6��@-�2�˘Bhb�e��t���I(��gb]�_�f+,�>��]�\�|�%Qn:���7m���B��?X��G��;hN4�m��r�?1t��V�W1a�Z	Qיw�cIϲ����b�)�8���D����ؙ�A,b�V[Y@x]�z�o7��`p���0ތe���H8�
$X2���9#Ű�����w�%�-B���`����?)�q��iW&��m9T+>�x&ϚuBڙO	�mC�����4�q�:?b��(>z�gI	�h^��O�V�1`"�jh�7��N����drDS�ՙ+�ui�SfuU�#Q��s���k3��[��T�ȢP�f(IyA���F9h`w�T2,�D> �u��H[9��8�F�؋��t� �|��/<`��� 
SLf3�����!J���q:�b�'�},g�T?/����Yf�bq�T�J����p�_s^;ϳ�n��gx^�3o0�ɍo�7v���\��m����m�u�;�L�L�L�x*:��fM��p� ���[Q�7]�"���ը�G����Ȥxzc�C��m�K�ٿ��4���]]�?n�d�m r���H��Hb��[/�P�����f����LX�g��N�hW�=�kTY���
{�oP��	���=i.�	3�c����&�B�B({�]�﫣�l5����0���3\A%6�(f(F3]=B���xul,��Q�����*�c86܂&`���J��q���L����`�]}��w�T��!}�Y����i�Z*�~��z���o���d����n)�_���&%��Y���\CU'א��`<���%��;7+TX)c7PYז����;�F׬�1.��A�����E0;V)Y�Ve�rI�Bx=�L��%�mu5D���7�_A^\�kW��(��Q��Li�	��N�r�N5�K\��AW��3���.zڨ�6ny����a>�>Q)F�h���~KRf��]�=��`�O���~�i��Г�)y�tiW���Vப����瀢"GSg��@���E(]a;0	Q_{|�L1Bu��>�����o����t����&�V-0;u���PG�2.��C���'�Ϧ��`�8�3��E����I��:pX�	�!�vџ;�T{�Z�{�2��k���[㛏�@���:ۜL�z�;���/�u3 a�Z������c�Զ���W+=M�IR�%w+�')Nfl����W��.c�X�5X�<��
vO�䞻�`Y)�C�j��A��
E�����*���(5��cL,'$�����^�T��J!�r��?�2�q�~/n����j�u����#�i���5����Z:�z:����KQzԨ�Jt�v��¥�ؖ!7lY����k�˼��F6Ԍ@�iDfDq���9d��I���°"_p�w���.=c�9nмP��R��ׂ*n�4t�h'U��,ir��b�9Խ+�e*��Wk��B� ��b97c�ٖ[�p��9���"f���#w#��B��L��gwH�ez`_��y��B}��h��9��
�w�*o*/���E��0��r�Ҿ�T�ew�ף{���0t<a���0cs}�^���kʘD2w��\[���L������T��	�x�)���ϩ�`�45Le�b��O�qj8�,%bd���x%�A/aϥ��Liu��W�~�R~�sC�5�����.�R��
`�އ�+�UXS\��U����2�H�H_���GrD�����nE=��
_Cկ*���w_���}k�5���vj�ME$θ�x(mp�U&]���X��
��W�Ӿۧ�L�e��m�_5�j�;
�I��2��#���.���1��}O�g�Jji?�-]��DE�����(qy.��`F�����L�
�^�u�\k�Jn3[3~u�9枱Z- r��O�	��s_�˕�=U�c��_�����	���s�׸a�O�!�20>�����t���/M[:�.x�����/{?�B������������wS#�)����5��(e+���Vl��^(�i�D�ɥ/�jd�RI�5-���u�_=�`3�TI3p_ټ��Kz�w�6���.�;�'d�Z�*S�5�o��.�y\�J�y#-�$��ٺ�z�2�Ʒ�L�Z����I��ۚK�??a��j����y
��m�?�����:x�!���-]c��p?r٩���^7��-;�A{
U"i���)M�!���Yp�Ԁ��~)��URl `���.%򵎼c~�RN�	��=�K�w�H�}������v��na�8�pZݩmGQs��PJ��@��;���$�R[�n���xh<d�J?_��1��K���^�T�
`�f��o�N��ҵ�q	�c�Ê#�ͻΌ��=��Oۍg�`�8�glqK�'��*s��n�/��ǧs��X�8��
�Xh�H�aA��`����$��z�o��P)>k'߉@��G�6i_�O�
Z�zI~@��k���� ��J�"=V�t4-���:�{�+9� ��R=>�,L��Bnx4#�s�Ŝ�e6���E���l�x M���E���c��������21�y1����%f�ܜ(� ��K
��	�k�-0���
 �4����l��{B����.�Ӽy�-��Jf� ��������RF�^F���Kc��H���l����������r��W��;��SȒ�z�W$��kżO�c�߫�/�w�/�s��jp�M�~B��j�����WR�{ WZ��]@ef�D�F}����Ӟ���ہPɺ��M�E�� .��y=�T�\/�#�#=�8�� e�Y8��4��$hK[�pp#�ޑ�Dg�i��}��)Pݨl򯭆][C�-�iUg�KlƖF���*>c��!�V)�pL����(���w�'��Mj���Y^k��O���0�P5@��:$R*���'#ڐ��/�@*Ӿ�`��0Yq�<���9�I���y�h�g�*��`Ŭ�֠������@��p�1�����N	��-6�b��\��%�ȕ�β����`�o9X�ti4�<�'�ElJdL�;o^�����Gܚ�;2�}y��Ϟb"Oj<�1@��5d��c��I�`[�^�ysi�3a����U��� ��� ��.�!\=���TE"X
{�~,���3[I��2g�V��n'R��<���F�?88p�*w7	M XK�UT�'��x5q��&sm��h�y��ʷ�!���*-2s�|���b����y�Q^���#s����Jy6���	2�y�L�9�hl��b�6R[�riBr�Q *
�����-0j(�����b�ESc�D�ld�e7Tf��O�Pu4m�㧋j��z5�eb�*���a�&S_�:@4�"ɚ.�F#�ma5�c4���xÓ���>�S�/��dI6�l�������[0�}.��_r����}.�ѵ��1읝=ȍ?`�H�sմ3�6f����P��$�j��č�e��Ђ ��PB*P��XImY�9W��K��iFC��h�Ja�{B�<9].��M��}��W���mnR��g��;��o���m�����;_��&{�������$�ܢ̥ߘ�wj�lj�nj�叟��S��d�3�����O'��&~�9���M]��u���
��Wt�{}?~m�#ОV�R�HҚ6Y��,h��w�]��8Z��5�r�����<��+'��X�%�o�)t(B!�V����gv�g�hB����./�+1}�5>� �ŚNMU��G��=?:C5D����vB���&dAl�H�M��/`��	���K�<�L�k[ٕ_���������'��¢�M3�PKժ��Vi����py7��X�(���%.�c� ��Pеv�9�٣G��*g9C����6� +�B�O���c�	GZ�[��vHZ���(�����Y�
n������	W^��\h������(tn)g{������}���7ub��/�kܼ0M��CK�H��p�Sh[R��23�/���o�Jۖ���#�2(�i�[w}[D�-5뾁���,u���1^�GU�3'�{)j"
H�
�y��������=��?�L2>]5�x�ª%:ٶ��}��?�l���w����Bi��wR���ɽ�����@s��&�lv^�վ�*�0�x��"+(&�g�T�Bt�EYy��u{���
~��|����`�q1�|f	T<�S]�7؇�2p[�c�ĐL���G�LH�b�R�ླྀ��
�G��]P)��&o{+X&8� B�G����}+��ܳ)�	?� ��k�i[��n+nC��{L��l={D؁\f{y�����ܞ4���_ׂi`\��p�-M��C���.j�^	��DG-?��` 9_Y����;FdZ���|��{!��	up��[�2k�*��9��画��,��2�҂l�N��j �'{�a��WC+>�^�F���]�v�|�}���X6���c=���)�Ѣ�Fl,�g����{s��Y�
���g*<���M^�	���B�#_	T�C+���A��І	<��"�U%Pߋt8�&3���)��@C��D�09#8�P�vV����v���}��2D-O�ߝ���P�|8q���h�t�̋��Ҫ�Aڟ���j<�PP�h�4����jD����� ���}��ҾM�[@�u<�+�<Lo'�������<�!4�Y
k?��F/���6ਆ�~���K
̑I\Q�W!����
��֍�A��\O�u��W��IN��B�vŽa�+uZi;'-�!��-Z��?����$��Um��Ju��E�6ԈX.�E	B� @�K|��oۍq��L4�乯���=	i��ϻ<�<���nwD�;S1[G
x����t��	~=[& �W��t12�� (J��x+/�c�"q����o(��x�#Fx�4�������B�d&`������';s�)�>:��N�m&R�Q��,Y�3��)�=�fk' ��ؑcN~!�7s0��d��P��k�x��#9;��[�Fb�;ёi��+���}�	����^���P��"� �����Z��L�R��4���a1_M_r��pw����Gp^�2�R>���u�8y��SN���mF��y[X4Es��-rGe?#��ʜӽ���C��K�n�L)�ΐ�D��eڿg����P�""�C�˾&���i�,���� ���j�;�!��ˠ�N�XK\��;y"�}Z��fT���䊪)��|��~1h[�d"���&�d����ͳ��:A��P��3�ˈ���WyI�����K�c�G�����QG��A�_��N��`?pyp��Y	�^.Z�C�Jg��#��N�[j��R�=�W��9�e����j���H���&W�B�#/+��e���?�'S�um�=��#����C�Q���x��0����>��b��,����_�2'y��4rB5�f�pG+�\��I1��|k� 
wv� R��ͬ��\m~�m�J^I�W�7#)s����r���W���,�]�hĎ�mK�����)"�����5?;��VI��ߒ��N]��=�<D�Q�]�s��,�#Fm�����c�1m����O~UYti�rlJi���ˡ�TR�T7�s~>�Vm8��E*�(/��w�f�NԵIj)��u�"�nB�-h�Fc���Z���*g&	j��胊s|���Te��~�tf"���|�}#��s}�|���z�,u��3�7�.Vډ9v�����g��C-]햘����4iK͙�ʖ.��m��Xi�U�����4^oU�bnj��2��&�q��2���uy�5��,N�~3I��Cs$�e�/�|���Z.�~�����՟AC�W�!�R�i)��=��c�?D�j(�������W���3n���|K����*�<��E������p�	��'� <�/26W�62 5�r���u#�͖�e���(�jΜ}*��ywq��3�.�f1��u����b�z�@XC*��{��2�b����Ʒ�B�(���E�ρWgN?��/h,V]�탶��FJ��^�a)꜄�:��h �2bd+�Qs.�Otf��F%/իۓ`�\w
�Xd�,��t O�7�H�vX�h�g�qf���Vg*��'�:�5�%&��(��T�Gsj4����kT�P����g�B��з,  WҪ p�\�%k�Dcҝ��*��rzS�H�)��%h�vt@�#�[{�����K���YQS|̢�N�8���b2�}��Tu�D]l>Y>P�ezX��>�K�n��H.���=Z0�c\]�/x;���,ר���>f��'?��	�׵1 �ڮ2S-�H8R�*\ >�K���Uz�q��KX�B��r�M+(��~aEB�\c��K�RTټ}j1e����EP�`.wyNw����!���TCx@
�!kY����`��8k���n#3�� �TF�s�ϴ�����'sa�=�یk��mD�R�d���P6�]4��{eǳ?$���uA[e~I��+{��_��pi]iQ�Cx�Q
��lլ�ɹ�ڱ
{ �3�$B���S�(&�w�q��t��:[��k�|������o�
�z�G6i~XV�l��4���fZ)Z��0��:��T�ζ�k�nI�d�8M�ъ4(/��?<�yg���̋�"6!�b���c���Ջ��X�?�g�| �S;u�%a4��ӓ��d���9|lG(��xv��֭E���B1��w3�Y���!2`�����T5}�G$�����@���w���1j|�6�B��@�%�h��6��K�6����,�Q�z�\�1�]����&�Y�5�41�r�}�=���59����오�EQ_	���i��
U׶�j�a}e�qxK�?�1�U�L`l@lu�KrK����Sk�`|=�v~��Z�:`��m�3�ZDZh�[����žf�����i:��������|�ثE�M��T ���S��W�-5�.�V���b��."C���n]h��9.b`h	�ʩ�/��F!D�ڄ�Tr��>wA����6��L8�Ò�AW��B4%�t�����{E�๼2�����w�ׄ���O�F���W�o8�x
�Sl1��2�8lG�&%L��rfw�n0$14|F.��#�QW�$�������d�ӥZ���)r��H�j�������Aw�)��r��c�s6X�c�5��@����,r�|
^ӗE�%m'��!�K:,�H�����g��ZL�6�RX���{;DNd�<2�v�Bi���gcE/���!����[rvV�@{��^ƍ:�L� b}��qZ�::=߾؏$�?;%TR�����sݗ3yzJ�:�$R-ai�fk����]8�"���Yo�`ҊN��*ӳ���=s�$��A����-
WE��(��V3��?S�O�Ȑ�8rh����u�wi`�'fZ���L��E�+�?����B�U���cu��;�����C`W��Q-ŠD��τ�3j��o4�۬�G���kw���L�� ��"In��'�x����ǺR�kS�sa�Bj���d����ߌ,������Az_�ɭ�T\��u��$0���E��x-�e�r����Ur܎��{R*�3W����XR���~��e��q=ކ:
cp@�r̥e�����N���ؗ��e��-��|Sڢ��
5ֲy\�@ v�@�J��ٸwⷸE��">�{���~?�0�G�2�P��	�nXnbE�mB!�!���j�d���e�:������+'��p��U*���U�O�5�vGP��!c.=���QsL{�y���yZ12E�ZA�A�t�:�1���	�jJ�,=��R�}^��!��l�T�K�|x� �\]��/��&�ig�di�ݷ��0��l���65�1���+��:T�q��tIw�؁��!L�j�^�tl�b�I>��R��0�A��FY��cǠ��k�Y+G��:A�O��?|݋���y�w����]�Ha��)�d������ �ꢱDM�ր�Rp�1�f8 �T�����ރG���/2j��MN��/�t�dZH&9Q������"`"�@�]�KyG���5��~zR��t����
�~g�H �4
[ҥ*\GK3�S���3�mU��.BW�($W��A�hS��KZ�����i9�%�C�p�Qa)2?�Ø��{�A���=����67�B�g���3�ډ�cbc��=�e�F������M�T�?r��n�Ɍ�eX���	�l$� �fgt��?P=A]�ٮ�+�	ىK�-�B�o.��fU�U��
=�^�{�B
�W���.��}~�g@@��j{�?����L�t�b��,#�}�R##ڞ�R���"�3fXz���n	�wC)�a��!4@����z��^��4��mO�:�M��Y��ͮ�c�aC���'�s���Lb����3���d��Cq�s���~}M�������^{�r�4-� �/���N�@az���6�h����5�������L�G����^\4�A?��ѷ�����L���)z�E�[D�~�~�y����y�h�QA@�!�G ,�.4����ǽR���Y���f}
�(�ȯ�#u�l+�	zլ���+�)Yz����{[�U�b=ߛo����Ee�J������a6j�^k�y�	p
����ڤC۟�3�mß I*��RR�+/f:Ġ��Z}`M�Rέ���f^��]Q�������X���OK�Ȕn�+�*����� ��ABt��u������鿢-��u��5�Aޅ�wB���JE���hg�����K#�jrhI��ӊ�N%�f�0��>��	���|�J�<��k��0s�Kb����',�,%�M��M��_�~}��v������f!Y1n̽�gص��Q��vI�W�VP%C��&`��<�9:y:�����ƞ�ڰ�l`���L�3���3�!�$dY=w*��.�@���dm��[��1X�T4��P���+/~��������;O-bL��>�o����VM��}�Kx����" �R�L�t�J�e���!iԦ�S�Z�~`(����2�9'����X�/��X,��^�^d��-��~C�,k���-��mj$n�����8�|H��-�I*�|={6�فnF�+h�"���J�%��҂#+���"��w����*�[<:��!�VE#[R�/���'���C��i��J��3.�L���Z��6��^$�hq��l��_@C��ʯ|d������&���Ĕ5xt�H]��_>˛�!W
sO�ۧ��Ȁ��?�Y�Ζ���GctM���M��'�;[`�� ΢�Z��Ñ.���!�^K�F��|u�y�`&z������r���p�S2�z/�o�M	��3
#�Ԫ-�J{��AE�)OL622�%|�����0i$���$�Pz�@���}���ޯW�^����BS��oT
�\�;{�����t`�Q��T@��i��yHL�����&��6��X���[���"8՟a�����<�_�$�$�Ѷ�'���[⒝�xq ��:��^�j��e���l�A�H�d4o�u�]ӄ��UI|d�q$״/��S{@��G &��'�@I���JG�7��c�6x雵�f5Vx�A��iDw��'y�iU���6J�+&���	�!\�O���B�]� �+�!M�4 ��
����g�5��m����աp��"bs�����ƶ1���
X�/	=6�A�Ү�����gF��z��6���Sa���S�R�	\�L��w���g���Gj�΃�1`.�@`~¬�����N���3�2�'9�e�h_SW�xa�I�U_] �V̝�;�K��"zI�D�yk�sJ����<��7>1��rG{-���5�rZ�U��a��7��a�%(�9f�䑬�UH'a�w��<7b�w��rN�C�fe����	:�Ux`Q�z��E	B�>1n�����O�;T��\H�ߺ��.�\�l3��j?3V[�[N�T�n�r;M�����:4�G��D2A�a�%��(����,�͕*�� PX$�犪��H|��J��6��i���:PG��]"��7���~��6j?sC��C�%*f�5���:W�`h�6�p��~���h�$�C~	��ܔ���S����E��)g�kI�R��˃9.|���=pLCJ�_��f5�iӸ\
+���R�����g:��4�q�E��\�*fN/�m�k���8��}q.c��i׃�5>�g���ĸ�Eᅜ��	��s�ٛ>��IL%��]�s�`�|NJm�����}�7����t��',~fjT��j��1��qˁ��/�A
�s��8�s`e�lDNЫ�~#|��}n<�;�:R��@	7�C�R��Y�W�������Pځ!�]D�G�%��Y�"�}���8elD֨ᆋO��;h��Z���m����@�حVxU՘�~'��YcDZ�_��B��  `Px�w�L��BH�� P�F��n���J�rdPz+��"t����!I��ZU� ƞ�Q�o��T�Օ�6�;��e:$����4����q��I�]�\�'sy�By�B��:i�]�a/�a���#�3k����i|`h~y}���v�	?I'[hbI�X����x{0׻:`m[cQ4m�\�2�	�Q��h����[g�t�Α�$�c)���_�ZC��-�v�*b��o���<�H��^�_ߙ��T��M�5U��f:���!�m݌_��ln�(�X��
P4�5x �I����j�&�2>�22'��i�ؙ�ҹ�#e��E��'�)���w�)��D�DE#u2�Y_��߅��J��2�]�'"(�U?wȜ9��Q�S�ޔ���7{�c�ô���2��l��1"�gw\am�'��[zY���Y)Wt�G�]�b�������+%'5�m,���n�w&w !�{g:Ig!O��?@AT붕lf��Y�+��T�Τ�?R��0�ͤ�CK�6Ӵy0��TH�%k�dM��RQ����Yq�>Χ�992S�a��b�c��#X2	%���`��$商G[LQ��.��\/4���C0Z	�*j�W� >	��jR�ю�7E<�����ͻ�K/9��H7XI|�e_T��V���gѺN
�\��>���P�������B�K��Y;I����_|�����Si,�a9""�例&����]��QIm�� ���ǺCgj,Q��D�T|Cމ��J���mXF��O[�S��i��l�O����	}̨��r�z!X�����l�Ψ��6�Xh�҆���hlM�3�'���C_ɋ�<��R��%��qt٬*u�3��dq�'�L�:�M�s�#��$����ua?	�;�����IE��
���pT�$#�O$L�����Re?�G�(B�D�a��oz���V�E����Q2b���tq�0f8���&��# ��*�[~`3m�K �
�A��Ti���K�����3p@�'�I5�-+��ݖZ��G>DĤM~��|�?��GW6Ez�G@�iW�o]�' bO��|=O����>��#��w�(5o�{�F�h1��]���"��s���(�����4<k9���6�`l�kc�Y2%�Ӕ��Ӳ*z*�M{\��t���^l|�_<�q2���ƫ᝗����'���I����\dW{��7��_���߮ �����WR��Jd��o�,�h*v����mؖч6�I������o�ʔ5pdGB�G>�K�������;X�K��K�F�Y��>{�Z���_���Z�K�����T�u+d�~ʄ<,*�>&�()��[�"Rb�p
]��=��ow��-���O��97�A��a�����˼�\��S�kqf���6H$����U�R����0,'���C��t(��p=Ѻ#�<��bye�x$��G��t]���X�]MYMJ$m�������"�!7�3���K�:�bi�5M�}5��oF��3�KB��E�^f�'�]D�UO�XNY������[=��ֱ�U/O�߃A��j���̣��c�������K(M�AÞ~�j�qF	��.�<�g|�SA���}uE���BHB�,�@���%����QGR���������9eRQ6�<{uc�����B�~n��:n�8�i��Ƚ3���ճ�Qn��Ǆ���p-��,�8$+=�ɨ�|�f��1�*�(����t����i����wG�Q�E�+����n�Z����|�f�Ԕ���F���˗P�6-�0��ÁaoնY��	��y%v^�����Gt��j�޶��qrA��3��y&@͗�{x��f������L{ܻR�/<up�A����I�x(ǈ/�U�̠)s���U���%�^[��|�t�~7��̾��B���譿�?2�﷋8 �n��I	� 8��{�|�(�ɿ�>�y�[>�@�T7��`��?^��?��e�ˤ�Ci�M7t6wO��,Ձ�_rev5�.�E<i���4��z��0��,��@����ss����HR��X;�?�
ٸ��	��ekl5cT��C���5��'�yU�`�}wr��!��h`�J�_W�鼧k�WTb�Ȓ�vŔ���7L��kU�i%[��
�_��r�V�)�4�� &Es�̤��)�Zy~\R���ԮMe��Vp��jJ�!�G��OqKLO�����/�rM�>g���.ґ��}a�"y,)R����`p�qG�B��i�D���Kշ�e���$W��]�;O�?B����`7՘Bb%X�0�!�@"���d��1��zuLww@[��.��E�S���T1:�?b�5�C�BX��p��Y���E�r���l�	^��!s�N����X����kз�Oo�ݥn/�����^c2��NP4���X�gp�@��^	<�����8�|�&z����l���96�S�4nK�FZ��]R��X����%���L��M9���}h��Z��͓Ky(�����D�c���+ ��7�ra~��,�V�	�)��!�e��]�\<�N>
�3���^\iԻ��a3��ÄE�����\�e?�TB����4�uz�n�iz~i-"��:������h/���`0�J�ͅ���,
���r?�P��"���mm��W.�D�i�z���<��u4I6��O 0� C}�J0�	|�;J(N`���}�E"߸�8�Q����	���ܟB�4�;���ua/�r�$OF�ը��
��✿�c*�T�~i��ji���Rε�.�,=��1�,��Rĺ�{lf*��/�̾D�2���a錃M��as���cM�:ըvR���� �$� v�X͵P,@�� $�`��:&d���{kx���II�㫀�(_!�	ѵ�s��9�p��q���l�P�[�Z�+��!Q�Z`;$�7;\�lifh _�q\J�9�r�+"��P�֤i�?'w~��7��^���#}3o��S��Q�8>���q��WH�I�S��k��?:�7������f����NA/�K@2���q&g����
	߷̔���ݎ����v�w�ڻ�-��H��}���4(ۉ+�〠K([u-=���4N�B!jL2%���7�Tk�n _C�6J�\(b��hCΦƛ� z|��	$��)a{���%�erz�#bn�g]N�H�dJY���)p��ʂ	\R��;�����@�Ȥ�$z�l{���S���l� �,gfrk�����pظ�~/	��	M�*�OH_��x���CW(���/c��ٔwI�@q ҋ&�}�'9x�`y&S��v��qS��p��\P���o!�8�:��A �R�b�o�3�ԇ4YW.*l�@Q�S�����{dr#���N�c�mj���=i{�����Ш��F.ZJ=��gz7��M�aݷ�������&�*�42�"�\��ܵ�_�u�jCe��vMS��
�|��ސ��qB�K-[5��u.b��M�{R,���1f�.뭩f���^���&} /���'���'{3k/�1�z2Lq[����5z��J~X�#���H�7���X��x��.��� =�<�~?z�WG�]���T$�������y��?WN��5,����Q�8�G:�ѹ��X��z�a�O�2`"#��%15�'�\c��gky��[p`c�=����w8�m��><?����q�k}W�����#*ۆ��LT^���0�"�;�V�{�<���?"�R��3t�����E��\% �HD� l��I��.�d1�t�6��ßM���_Kd�CډX�����&U<���y?�n]��PV>�eƩ�|Hx��8�(	��͐m=����`m���u>�;�+F,R����q�=��!� �IT�џ��U����t�/pI�tM��q@�٪��h�ǎ,z2]�����{t�����@��D��^N��-D��#s��������O��3�n�%��z���>ԪM�N�}�㒖W�)��̒)R�a��G�H���fN��*���~��!��s�ѭ���D'H��l�zMh�+q�<����p/E�M�l<}՜(h{;C9�p'ȋ|A+$� ��ɑ���c �ĸ
r�4��yhyeb���w�|]'��W�o��p�߷9H� R����O�lq�j�gT�V��iY�Ae?ا ��e��\�A�����Os�,U�X�\����6� ��OSԖ''��Խ���@�K������;e�������zx�,�oRe��Y���<�-q!�:9ן,l�Ie�r7�Z�?�L㻠�%u��S�����5��@�Վ�	!�]s�1�G[��t������>Qj�E���G�w2J¤e5��3�k�"or����0����|A-]�H��Fp+.�PrT:�౵;����Y�c��F����C3ߨ{)��*���3�T��:�>/�
��^�q�����[¾��,׊)�k���Cr���8Iz���8��chX�o�<ʝJ�G��+�i�GA�eÄ́�H���%�3�{ R�Iw�ȒO�ߟ���^��s�c�&I	ɉ�K�!c���Q#dI�8//n��`�� �pad��.�n�1��y� =Q�����e��g�3�����!�^�R?�+���r[�2�u���-��!/m���M��Y���:[�3���&Z��Ho:C�w \�ep@r�`'8/��}G@�3�[ԝ_��wU}�iњ�U@K%��H��2�6Sײ6�HI���I��"�	p�W]��JHt�7i�_�$$:b��0���S��y^>Dl�7}>��438�#	��e�IgMTHyޟ�+8W���%�N���2Q���e2�	�F��L�3*�!z>g?	�c��к�`�ob�/�P?�O���4�nIy��y�:�Ţ����W8�����o@l�H�� ۆle#�����Y��*�OW�Q�)������e�F�P{OQ����ĩm��F�d%�I�w���A6w؈�/B�y��Np��`~	^nH۽i����k�ܱ]���8����0~����=M��r���(g>\�@��L�ڥ��Fr�~&�*B=���|��X;�G�Cs�Cxzj	qF����TV�T&��w����=���^��i�D�bj��I�Ce${뒝m��P���鄦�(ۗ�mD�*DU=���V<�;���1d���繳A��f�2#�q�Ĳ[$j��Ђ#�
�6
A	ڝ"�qT{��7'f�9�n�{��C� �"�O�%t�"��&L�7�2t����샤�*#˰�)�L�ԩ2�Ҕ��-٥�C��KO�&������ba��o�Vs��m��S�ˀ+���t���h �}�Y�A���l)�LoZ$��p���y�h�aҺ�$[���8me"nO^�C���Ӑ���1�)v��ft��`�\�A�p,�������W�/0���|�d�<?Z�Dv�BJj�D����}�S%�,�x?�r�f�`U�@��������|D�#
Q�:30�荐c���=
��}�eN겣mLɒX�9<է�xx��p�r5���N8m�)���M��PDSի��S̳?;�[�)�7+�1x�jJ����v6�L3�g�v�_W�4�p`o����R��:�[x��N���(�٨�U�q��� e����T`�U�y��L��?�B�b����p{������O�>�����B��='(<d�^�!��{lм�(5�p����󜞢���N�m6�V��\>z� ��5�=��������̩�\�R������R:P�ց�,�L!�d��H�B���s��^�� �9}��P5��,s�i�MV#�=��JSo�Pog�F6���@����z������LE3�<S��N���9����+p��v���T--@��K�I=z�	�Gč�R��dز��+�B!��f���ӄg��uKi�)�w�*v�T+�vQu<�!+�s�3�X��r�9���_�&:c�F �V�?�0�0n�ohV��jH�,F��7l��G�i���W;,�E��Qm�1��)�%ӧe�J�I���T�������a丈����������H�Nl��Jp�s�,I����|�I�n�g��%eض�w��w�7���hdZ�V�vE9ih�T���S7q�]rT��tB�Kh��2䗡���nT��+��<�@z܅�C��&�{P��n�1�� ���b?�:�n�u�? 1��O�f��&��2)�T�+�U<��y��3b����_2�T��6�׽���AP�Z�@�?�|�,���/R+�G�m�Td�>��V��lM6&�g�=�_����ǧ�af��f��9��߉9�vW�5dZ���+�q��es�x{ ���/M�zb�8�����\�d5*�J�t�b6~���ikO�D�#�s����#���ߑ>�x�'f(n|�m_�6��zYĕ���ph���Q:��6W�����F[�~�`��J
�t1�ۉb�s��8��2�Kw �ZŌh�YS�1��EeƁ#�&rjN+sc ���ҩ�����X6`��y�Η=,A�6�z����j���w�c=v�+����7�3eӄ;8{�ץ�r⁨I�7�X���ԉ���>�3����^w������ۙ�>[�2),�AU���#Ǚ���S�������2%����4���ߥC�~���
��JÝ{��M��`U�?���T�N�C��L/g��k�ed!v��6���� j복��7o=���}��y���*��rDe[0�H�3t�:��֮��Wz������)3���k	�Eᓮ��o�W9�	r�0�?Ӄ�ں�3�X����;��A�b�*R�����r��D�M���y�}��@%=j�7CBW  ���J�9om��Qќl9��^ߎ��w����J���a~��3��gN�¡�-v�Rc:��c3�U���n��1��bi��r��g���8 |I��S3Wy*ΐ���$u\�������-��"����z�<�����? 5?0g�+�7�a�v"�w���R˙�}D8��R��{�V������u���7����e�skԍ"4^Q�q�=�e/�/P�rY���&�']�<&�]oW3F{���)�7(B�$�cz��@�S�|��3{��Y+��D�#�P��q`0�����w��֯VB��E�M���li�Bh=Y��(���$%�xj�5�A�'�����~'����ʧ��8� �5w2)b��5Ya��V��e����Q ��M;B�^�4�Vʢ��67«�t�j��~�4�~^zǢ�������h��:0��O�� �u|G+�Zޖ��Xk+)3�:�������܂�ȁ����ʔ�3w��V���8H`Ps#�-��\Ё��?�`>g�Zj�;YRN2����ׇ�����c��z��յ��f�xEr��>4�B����
!i�^�Z���[�3�+��(�zB�&��`5ofK�/. [E�>=�u��0��"��������´��F������k��T^ �K����˟�lp��
� }\���Q1�?�t%XQcC��*�/M���]/,䭢phl��ɽ��C�\��MQ�a����q<UR�G���I�/���Y`�'	!Il9"���L[����pi�(ގz��ň���w�N�����k7� ���"5�S���ڭ�n�̞��HvS�����U�W�6Ze�j|��K�x�o���"W|td*uõ����$7���6��Q���#��b������NB��bpЇ��ŪH.�~�KG�vQ��PS�H⠎&w#\�Dik:�T�Y�,Ȍ�<���K����ѣw�#��W�̒�,ښ+��,͇pcz�b��O������a���Ni7��s'j������dB�b/����2,���D�Tf!��.	š�5���/z�L�� r4�ޚ�X{q�9W��<*�R9��{���m7�վ�#Wk�"�gA尿��v��+"������dQ\�Ǹ^��!h����a�:�(<���鸰;W��9��脃&��a��Cv�W?sÊ�,�QJ�{;�����%ڬ9�AK�ơp�g��S�1>����/������mf���������SF%t�b�	�'3`�2G]�i�
AV��w$�)��.ec+��x&I�Z�k ��^t�����t]EѸ�����ۈAEd�g�>tXj�7�O�V)+T��5	���@���Δ#�M������ l�1��r��И�� ���$������	�ӭ��<���>[fj2M�e���$��L�Y�2�yRG� f�/َ����e�,��z��?�0�%��	u_�
��3�/QxC��2Z�b-&���1�XR~���zy��gi��\��2~	�|8��W9�m.��`�$&��5Բ��X��~=���?��qCCC��'�90Bm'�!"
 �'.�SjR[
�Ѷ"�$uk�6j��B�o��)�{��/��+�A?;�~P<���&�k+�Ӏ�RIE�E�Ė�ɑ��%]�f8�;Y�L�\�T��N��I���:vLS�u�fh֭���aZ1o��y��?����M��0�1�&z{S�ErpdT�x=��B8R�&�o[�/��KE?����YLc#5���Ư,�]U�^�������9��-��=j��}�����o��� `�F�?���Eߎ��> ��o�h��ZȯױB�n[�0���!��"�iU
G}!�9��^��-y��=�����P}F����2id�X�u���QF���;]���������+��ٱ_��^�����F*��5bNV�6ƈnE��;��O��a��Xiq�+����$+��b��i�dó>��L��5ύz��Xؗ�� ���Dˆq��(�"^���F M�R}=�bʿ_��m�V��!'�(X3�"5-fFy�MiN�r�� ,���6�Rp@hU8P@3Ú?{��ɪ�F�tTm+Ɋ�[�g;�)���=��g-~�d��ej�l���[��;�X�9�;�Ȗ�@o@�|P<j���� x�@)֍��9�*��L��]��"8�y���E�� '(�;�,?��M2��?lK��,��9��Gſ�ʉ�Cc.��p�!.��T�O��oA�ql_�Dg��M�.ɷ�@+P��v����G�g��E���_�&��Z0�Û�uiα�\G"d�(��Z=B^1�޸k��@�H��N(�m ���:���0��c�Z�\�*��x:v�[D%�A%���1�����ʉ�D���*&!�đ��7U�-�2�y&aK=>o��D$���7Ҏ >rJ��8Fm�"��3� �QZ��}�gr�q�¢��:�/�;N.2�
�Л�c���!�/�#u��ϩR]�%l�t�`���ݥ����#�4M�i==í�}Ю�d*�N��q
9Z���v�|���X�qr�ש=���M���ʬ��Ax�#!:#E��H��6����B�~jE�g�']�u�|��)�.g{���l�z�_�HZ�2\�G�DGM�F���Z�h�6]{d��\�W�0Y�)��sH(	���̨�+�N����{��z_�,0f2ga�����-?o6��s]��@�EA���2/�R�\o��Z@��=Ԩ����*j�ܘo��O��~��[�ѓK.<.q\�v���H�~���*��ѯ��oo���vy���7\���+��eԄ���g;�ð�RF@�ͅô��l������A$*�Q#ķTp���!XZL���@���0�^gc�wbJ�x�&�A�UUmAJ��:�D��'�V��,Ǭ-��~8���1��^~��f�I��(�g�� '�*���t�<ŔU�*�����`�(����0n���ϵ��\�xPjZ��Qs���(/|:�rq�#���.��M���c�UB��YbUg2ё���E�DJ�ԝ8[�ydO�N��c�v��E��f��x@bYJ�Em��� �ƻ�Xt_%4c@J�	���3*0���lQF?�t�N���TqZUD���DV��;I+n�$�Bs<;9�2!&q�5�jFt.rW�<�*I��q����..
1�d��DXJ�����Q�� 4��JJ'L=ؿ�gFy�ߵt��7:���D�JCI��9�זK�25�x$���V��K�~j7\�q�5`nmf`�`�K��o4Ո}ߐѕJ���M�9h�s�<��/��Y}M^�is��y�+x�J����BAz�ϐ�h��h�"�r�.Nwn�/��;������Eč[.:Yj�5�l�b�m�5262�X�� �<��5�ML?�9���cQ��@u�/=��:���9�0<�j�;v`�eR� �1��3c�z��|���%�tn�Ф���[�
[
%�b�T����������{vR2�&��!5=�6��[J8	���}�5ْ<�X�s���k !Wx���/�cw�hюi��NR�Ғ�|s�#�F��>�������W�re�؈M���-y8N~�q���Ǚ{I��xj�mzI� ��0�����d3������:e�m<GWY�"�lܦ��*B����t�91�56�	1)����94��%/!>F���k�V�C���i�9��>�O����z'�C�7!�Fgީ����F�E%�lnc&�FOv̛"<O7�G�_�^�m,�ћ3}�㋥�G�0��#;�+�=BL��B?�����ʮ��Y<��l��2��� �RX��^d+����b@1Z���$�?~P<��J��&�!+�f7�<R*s�(������+�>���ڤ����whv1o�:t(gc�!]4��LM�4-����-D�X���������z����$]�>7�-���,�ϩaL:�&D�&ǆ�t�|�GO���l�p��ߵ��]���9��-�$�c��zGl��c�V�A��Z��?�w��4h&e�����Ӷ���y5R@���gj%Y,0KÁV�{h���?��������녥��K;!��#�򤀳����+��7Y-���>�yԔַ�`����*��I ���z�h�OM)�o�h���9�U�IBd	���7���L��H32�PW�-���ɼ�@)ÄT ��Yvr�,0g��+��Qe_���k��!��J=�k��Z�q&T�]���ۆ�Պ�JK#����yH+G��5߽�s��F[f���?�*�
�R��ȑ>iR���ø�}�]XڋC�H��!�9d懂<��)���^~d4 �fQ?��F�F�Z;�DM� �m��,�l���A�ȓ_�ˣ]�$9�`�Z�����a/��������-��������+^�#�)�Q��&���T��W�r�����sr~f�h/-&�6���`��|�9M��wF���0�0�6Ϟ�4b����P1g�tP����4�B7c&GM��z��dԕ�t��QQ8�/�uhq:Ǖ�5�4ܮ���M��	�U��z�ީ͗m����_w�c}�đjс�P-���P�ݽU>��p8ioВ=�0���\&9���:��JC_z�X�sis
ڿ�P�4�M�+��n�!۱�I4�{�W�s�Q�� ���d��"ٳ�����D��p��u�S+q��{�3˷[�EjTܨ��tʚ�oӯ�$���9|�'�Y9��Ap3�Jc=cϛ����E�KIj;�G�e#w�
ӑ��7Q�`mwK��0����9�:�#ɎOlz������٠�A\u�7�NW <��������&�1fQR�}�/f���g��RK��l��][e��0oBXv��{z�f��HO����ܻ������y� ���ҽ�ڋ�M�3�r�s�ցP�/w"v�wsq^w�e���ͅ��ONwev��*0Yt��<�<�b( ���^K6�l�(�)҅���(@|5~3i�����F(�Y���:���y�MJ���S1�����Q��֕�p�<u!�s�|<�aeh䬨��и�J�~׹��H�B��a,��K���hV9k���8c(N�Ɩn��KR�1T��p�|��)r���=<`��N�BV�@y�.}Qp��k�>�=�S-����������4Q5�x�O�VE���iw����E��u��&N��Ge��J��gkg��W?R�`Eo�o��	a������˭�WQ0���5x�+n6>��IE��]E�����q�FA��-y��ec}lNF`A7�d��5�^7Y�ig�`	��V#�J�./39��1��]���|4X��@�
��J�5�N�~Gf]Ë���c���� ��������
� hs����������C�ڧ���Ŭf���Tb�����>�R��P;�xW8���|*�oc���`(��0�w��'�����_D�876>Ȝ,�z+�&�;,[������5X�?�XC�Կ��/*4:{ө.�+�	ڟ'@L��f�2�l|�Ư|Pf=��B�f�WG�b쾍$Y���'���J�P�z�4���RA���iH^����ʁ���+%�Y��lI��	-V7�)��C��x�Xޙy�KmN���nP�O�B����JfH3: �7[b��q���eK�C-��U�����cbx�ُ\�~�w�!ܛ1��=rϮ��A���-�����f ��Y�] Ul���ob�8]V��wކ^�Og9�/�v>�}�(*q�ի�.�V�
9��N<J�.]q�3nhq�t��[xd�{�PN�)8��L�B�����,��Jc���%o�S�/15�����K���w1� �_��Z����J���-=��K�'�~�k?Y;-C'�����ђ���;	�?�P*3��~�n!q��n���7����34 '�(jN+)��љ�N#8:s Q	���ۥ����DNf��,�8$���F��nɱ� ��diU�����]�8���ԧz�.٩:- `�X��{Ü3�{��2��lT+�	"�p�u�
E�nQ��\�����L��h�3h��<W?�͎��
�j��u�w��Sv�$�O�dU��ǌ�Qœ�j5���K@�\	�0�=���f��'R�q�iz���|��3@Z�m�����������h9Sl,E5g��g�9(�����tl�E}�j���ӷ�U�mq���W�=	&���.v�|'�w�5f�.�h]+��p��H`E�A�>s��������j�j%�~�#r^�	�5���v�����{t��"�8�V�4$���3<�x��z2q����vS�,���3�x�0Rx�S���KkT��|���>iiV&t�s���tf�E*�����A�j攠��3��D}?ơ��]oWh��3N;Y��Ʒf�!F��}���Г��Z��T7�rkө�;M�nU�_�o��rNf)�չ��Lxبa���g�`�Z��)5����K=blr?W:Ƴ��_�x��C���A�J�+��۽����������*?M}�g��� ��ߊ�P3/9c���i̩�+r!c�B�]�r�b��=
|�$��!����:Û�d7g�b�<���Ӊ5fBE��_���ƈ�DY �s��O�*߱��	���V�_���X27� �}�-������q���Ji����ܕ�=�#�׀0Y�n����]�a��Q�W6�t�J� ��"�B�(F�����)��[�w{0;`���>��ʛ���AX�3Q�X�yʡ�1� ����%.ͣ������ wS�r��M��f�T�b�w�ܾ�, ��xɗt4� }��z�28R�\�^�X?k����mQ��I�h�� 9/���:��������>��f ;�Z|��	�M�-�`K_�G�� ��C����|o�1�zr@���(� d�b�l��Y��>�+�D�f+W��g�k�o���8�E���B��Dv�\��"SY��)��8�	[po>�(u���%�o��{�V��G&���ʳ�Ǫ�X �͈T�W�0��jEj4�Q7bP����1��ѐ\5���^]�qv���AI	-t$"��^�ʽ�Ã��6 u��H���Q-/U��<r�D�d�uk1��7��������^��Q��s�L�����L�[��$�#k%B�Ѿ��R��m�FL� >��7SrH�67���� w�A��x���'�>Ü��/����-���ly� KD��G�p��ʶ��-VB|b���G[2Gg�a��Ԛ��G;с�K��4	��=0@�\b܏�<���P��.�kCX�AP����Ě$�9�-���	v�Ԡ>^��ڸq� }�/Wε�
س�޸�0�a�U�7�7�4Q�V-���m �Lqt�MH��3�r$)�+�����wD���]��l_�5l�3#��v�݁-}��z䙞5x�6�&��O���Ǖ&?�-e&��sA�B����ʩ��_��׌�}`��7ڟ�b�R�e��(��\ܻ�H�$Yq�Od���A|����l�%�ǆUuRØ�`��T���>�o��N�4��W�[� C�#v_y\�;��b���$�����ǯN�S)㕪}�-��������5�O���O������CS�I6��EO��V�EcE^74�����)�4�E�Xڤ��z��4?K����������h�����04�F�=K����XT}b���Hʟq��f�ŚR�� #����K�GǇZE������&��������������#�F/�AbfJe3����oD�����ņ�e�y��}z���5��hw���ߜ鷔;�(E�3�g�,�8���>����AB`8��B��5p�|����~_�T��cI�sDr�ޗ�}�8J�'$�����th�����qOg?�m�����>*��&�}v*T2��|�g�ׯ�s��q�3p�b<9��0?V~gM�q/��J)<�m����$�9~Wn:���M��+��k����1@P��]�=:�`(�v[o�ET�z?yI�= �����Z�%rK��$���Y�x�S���2����O��ƓI=�!��&0�^=��������t/v�N��X=�^�q���n�M�!�1v>��Q���s����(�NݑS����x�	�QK慓����X�_Ba��Î@{��b�4aI1��	K�ڌk��d���I`=v'y��������*���9�k��D�v�!��q ��R_�-FKIЧ&o �Z���!��}���*e�:w>��ʎ�c��J�KA~i��7/+7T��PTX��܌7�	�6�0��x{�Y�'�$�P�P���~��0&�S���γ��F|\n@|s�4��ryc�)�
�n RG����W�Q���pl��wӴ����|uUJ�
�OӲ|dK/��	(��L�IO��!�K�h���!�W���`�z�rG%� ���Þ�<D_�/.��3�*}�o1'9��K	�ł��:|���;	!T߂�[�_�\+��WƎ�^����l���J����g 3�"⸿jk�Gfwt��/�v#e��j]��� =�O�s��n�T8�o�rF%��U�����t �$.�+"G1T\10+,
�V���p�	������=��9-2V9�p�.`�� \��=�Vi�`�l�I�P�B0��p:EB�go|5�'����%�/�~��)�VW��DQ�6�-���X�(Կ�Q�r%��|,��x���JG�����Tκ�Arh���̈́���-3�b O���32��"�J�1k��N3t���-� �G(�ٱ�0���[��i�Wk���}0�JZ�����uͭ/v��N��]@��선A����Zs_.7ۛ��.a�!m�vr;?�O���}���ߥW�}N%�C��נ�5�4��&u|Ǆ�ycc�7��d���2.�
Z�h%]ޠ�e�߽�SVʱ"��H���	�"�F�o��Ӳ���/;b^�m{*/�s	m�Δ"�ҏQ�5����̐��޾�g�h�o��pcbg�U��}ߗˬ��v�j�pKk�TO×^0:�!/�&��Q�S�>՛KI���aЩY�C
F\�t�{�ٱ�'����)�|�o15�2]u������Z��<iUa���ϫ��xC��efv�9���k����#G�4�2�n��5��9��>�����%X�ǂ}X�g($��p� K�:�բ�=����|W*;clV)�j@�1�S�z�����O0�^Br?x�3��E��rJ�AN�&	��̌f.N�wz�V5u>�X�s������$�8�6x$5�[	AT������`���ƦF��
�n��<��<�y$<����_@���ȟ���_~X��A������=�4:c�FՐB茔�Ŝ���Ƴ�M�R6^T��k�=�nrqh�nh����$$QW�N����@ϗϙ1:Jϔ$z�~�x���e�H��ހv��m>x�j|��RtQ똏o�a*G��|�5�8d���7��斧�������Fb��s���Q�"�r�k�eDS{�����L�E��k��7Ao֠���fT�R֜C�uEN'��V5���G��>�L�r^�c)*�@�c��I�O֊w��/`6Y�����F)v�@X���4k�~�������>f�_&ԇ�vRL�|�{��8��L�^��?z�����8�Y��KQ�x�^�X#ΐ��x��Q$�ZSþڶ�����B��U��~-E�-!8Ddh�N׶m��l.��@m�r[*д�Q|&��JnP���w�h�Wnz¨"Y�����W��	O^"���*v	w3�~�B��33�:�;��ܟ��Lꐦ:���T=u���0�X�Q��ӻw(������cai���i��j;vM�Ku;j`��H��^>����s@��_7�d5�����٪y�h��Ɛ�gd(T��|߱W�stxV�P�M��:�ɜO�eT�폙 W�Ɔ�ئ��dJ��=c_�N]eY�B��q�A�V��v9X)+�q~b�N�9��G3����<!��>�Z=P�+��~�3dРW��7�^�/nwų:O�h�ѝ����'v�a�ch2�a�+&��P؝D1�H��"H��J��\6�:C��> }�~�wv����ob�-��<���i2�-Y�_���E���th$�$*ug@&wt�z5a����VAMҪJ�������j��5%��ϛ����W`�ދ�E�W����cRr&��+��1��ӈ�g}~�F'tI�k+��ѵ��54�|�����y����-�IHw%��������n���]����YT�?߄z]�$�m������܀���\q�f?��5��2m���]�W����H;)+�:#��IPc�7��zw;-�I4�������-�UvF�	��!On�q���`x��e�'
�$���ѭ��j���z�|jH'1���5��3I1�\��%,������t�(����	��v�u�Z&������tF�=�?����y�����J�"�aD_������9H���5���G�����xc�j-�2T��a�K���{�g�A�E	;��o�ݗn�j�� Z�*�Ė���OfT�4�S�����$ڕփ��y���)A�o&;��[|��37'���e�ݏ�mf�dA��@��������G��l���Eך�[_[����Q��k��D��%�	�@H�;=B�����T�
Ya�X����E���,�#��~LY�����Qn�(�!�7�+wR�-b4u��J&�ݎ<%ڤ���j���鎷�O<�D����OQ�r]#�~��EŦ{| �i�M��"!��P�>s�)B5�ύO�j��0�
��#��/�p~��0\E�wDޠq�3���P�r*�<6bD#{�90���`++f���?�����%�_�ď��@�w�.�o�ik�[Ƀ�L9s���M([���f�$lȱҙ�h��F�t?IO��j�w��%�5�:]pn����	R�������fZR4�q�42~��RNš�h.���z�S��f��4�ma�Σ�B�`�,jY1$z0|-U��	�w& �Ϸ]�cU ���� ͹�/�Ed�}.Qʊ"O�;؋���&R��m�F [4}��io�G#?��-��z,%�˄<���y��n�%̘-��P�k��⧛����!��/���;�����|��`��M�kKT��;af���t:Z;��}��u8�g��Ā�<���LT����!ћl>u�(�2��(��7�"&�܁_F}�#*HYF~��1�ݸ;���bX����oY��i�n�XIjk�#+oM�ۛdҿS-;����{�!$�n1��`��5������V�=L��6y!���$����G"��݉p[w�̏)2�`[P�ҿ���K����s���n�w��4���Zu�&s.�j�{�	��Nԉ�z�}��5�`��ߣ��d�$5�y��z�j�ti�Cns�GM8����;?臷"�7�I�rz`巟�Sg����%�1s{?���E�F���5S2��VN脻�G1W��_ lB�sY�@~�^��y��g&��yU`
�ы�cR�~kN���%NܐK��pk�LU���;�����ֆ��%����n�� iā�������V��O��ѻh�o���V�	���A#�w���)��>����0��24���`�q�-�&[�<+�r�LJ,�>�wM����/�9�'t퀳��ϒ��լ�;2:��[jr<I��ݎ�2^@Sk��8�=Ö&�R����t�5e'�_3�3w|tޗi=�^jB�=����)��~���{-n\�.���+� ��	�d	�pò���8�󙯿� ��R�s	5�=]�X��+�]4�1��w7�)�fpd]9dJMẾ��.�4Y�Q�h�h���-"2��8�����X �[���::�r�虙��=���A!Y�Q���v`��t:���	LO�x�2}躉jF������!*�{��`�ڇ����"ƅ����M|v�����AWu����	�PYA�Υ�x�H�4�A��&����:�U��|M�v�"�����22�C#U#c�S#��F�ڌ,�~q����F�1�E�j�P��v��1��/@�T�S��^��V>J4;+��~��7���FV��~������̢��
������­�Hw�i�,>��#JS/D`ۦ��
 ���[$$w�Ă=mt8x[F܂�H?�B�s���ȅ�{��Z�:���K*��Ii���p߁�z���+��싑�����{N�@�/��B�����z�>��l�掓?�h�:�nd��|��f�??N$����D�5,��T@,$�L#��F�����X��&�}B��!B�A�	�	V�y����(��ꈇ� ���$ָͰ������՛e�mW �����A��l�F�2�@��/����
���O�~Z�Y��~��ײ�o���4{��)��ʛ��~�h&�D�]�Y�;�'� V	�隗!(�y���djr<g �����I��tg,0	RE����,0c��}Vٚ�4^1�f�V�قmh[�d�)K)Gѭ���e��9ׅ+b��܌n��d�ǃ�0W_�
 �.�5���X%x�p
�ק_k���v�T=@}2È�I��k��:A��U��^2HP5R����I��q<��")�hы�@���
�Y�5���v����ͩO�0ד��������I����/��d9��Z�c���+8���1a�����9���n�`�y����ۂ3O�[N�NK�qg��L@@s+Z�,�b�J���p�~e X��0Д=�Bg���#�t����7���y����$I>:�l�"5��S,޾Xi�#]k�;H4/�	f�mRK��w#�&~���=#ga��;v*���:�|��ݠ�P�������O��]�
�U5��'�~č����2͇�]|�s����y�
����������w����c��xj>��蔪MIZ�QQ�����h�&�5#�ńM�K�v�Kc���t�g��X#}mVy2�#3�W�RuX:��/ﵜ���L�T5�cˆ�0r�0�~� n�����5nU2(<-�s���+�n+�������+���`<���Yڿ��|�*��\te�k{��#�%ş^��������'�8I����|��j?��/j�;]�*��8��7��O3�=�>��~2>d�>���B�<r.��lZ�c〮�#�>Tf���5��W��2D�.K�W��h���K��!C�r�AE�FC���ە�|D�2
 K���[�|x�ܩ���i���<]�>�a�-��[����սY'�5��I�L���<B뭇I��0�����5S٪u��m]��B�>S�����O��}�;pa<� ��\@���j[��R�FĞ��z�D�P�e�P��(��� Gl,?��+}5��/��jM4)�,ʹ���i�xA�:L��lK	#+]^r�]n�kxo!~{��f��������Ŭ*��"S9\XӖ_�/��}�0�I��]��ֈBL�p�D�] F�F��zyM��7N�'��16��7o�����D������~���K�i�x\/�v+U�Z2S<uRqq�*C��1��Z
<���HǕ�S<vØ<�"m�U�E����$͎�Ff���q������}q])��l�V�zTB�ɞB�6�d>/"Cx�u^�&~�쿃��a�8%��p�&�������,�`��9����$��`'����:�9r�I���e�����(��둚�����֦������>�mT;�4G^4x&|cv��ZZ�M���u��˿`ق~ IyG�ǟ�m���
�<=!7���+�[$�b¢����9o��H��^NJ�U�7�=���E�cG�@"�
��WYW��ք��YRc��eVN�D�7���� � ����u�!�f4��qX�Fix��jC�#QBy�2'���c]g6��/7�������r��8.B�N���O*@Ì�([�2E�&ύŀ������Zb_@�,�w���R�:	�Cf��g(?�iZ֡��JM?A��%��9�О�ld�8�����g�v�����Q ��~�6j�����4[��k�*���� ���!D�:�e��5
 729�\=R*I��񔄔�D���팬��� odR2�e����qZ�|%�\@�rK�O� �o�i�~Y�%�/gڋ?&A�������I+�G��l�*}�|������kgS�� W��9��dV�w��ձ�w.���!\��1N�H3p{Xf����2������Sv���'si�mk�:F@��u�i��W�.�zTe;�uh�_�*���?=����CE�5L^�����ui/�)Q��-�w�6�~q�����;ރJ��B^i�u�q��O�NZw�1��n+�������?T��z��ӏ�A�o��-�:�]������սi֗��͕i\�3ԙ��'
��I�v��(~��^���`�=�5/���n���;Ts�jsuɪ!��I5����omÇQb�z*��9�#X���ڂ�8k��6�c��%�IGrûy�\���W���p:oSF�
�����d4[#(G��7�V�Q:6Wy�V�E,�SY�Y؊@���Ƅ?�Í�\#�s^����0��F�^�t'��D)��MR��S�����'��Vz�N���>��ZJ�QQ����л:X*��<p>!��-*�f�f��|��K��~�)����7�>�Ֆ���9M��B)���vV�.�b��[��}|<x��ݢ������h�
˼Uf��D!-3�<��X���a�ck.�:N��~\gw)M�g�C-�T�J?e:�?�k/�A��y(4��#�W���a9��R�!�mU���:��oL�I���8�9msg��(h��g�o���u�5��/5}K�dN[E�f��^��*`hQ�d<��X�>ȯ�V�p�$f�=�ذ]WP*�;��"$X����@��ĜI��$𬛙0�+E��)���-��.~�F��'iך'ԺZ�4G��טF�;��'h+�oU����}�&=���%o���zbW�q��y��, -��y_J���}[�A��W�O��g���@E��!\��	v�Y\�,�j��-f�;0ƯF�Ɗ<r	op�W�ql��hZ���e���'���\�b!yhx�$Q��.K���S�W/���X�'�y���pg7�͔�r4o��x��8��i(q�7C�]ȳ�jWo�$i��.&[��dD~�h8��(t���4�K������ãw��]�y��NI/(ą�ޘ"$	��_���	�m�!I�"y�&�%��g�pT�[d�Z�~���snI?��N�/�F�����k�P1�#�hR�Q ��$�P�6�r(��^�5E_�3����JGB���ۧ�u�^�3���d�����hP��9>����{^_���t�@�"F��	���E�b��:O�$R�v��S��J<��mMm�(��O����?ɩ4�[�'�LJ�f�S��������9\>���pk�����9�ϧ���6��,���,.*�2;�ϹP�"�Ks\�������p{q!z���A���L�Y�S����B���w�9�U�I!u��`ĩ�@���"��������6-�5�xc02{ӻ��'�b�<����JM}R+~��$�77�Rj��wKKH�ݓ����⽔�Ky��c��}ƽ��y��RByU+Q�At��n�����p�Q7C����٨�3.\M���:�����&bX���MEh����uQ� �<�R���g��'����^6��!`i�{2�s�;t��.�<�խ�������4N����u������=��PV/-��r��Vu�p胐��Q�7�wҺ\1�Ƹ��c�G)��-�'!�+�|y\
2uMG�7��G��O&�M��/����i*����ڼ�s��Ux� ��9�;�ok��!��.���6[JJ�7_�4IV�� 4�"m�ad� >���+�N(���f�7%��2;��.���rŲ�I�a�9Yz���[֯�C��ɐ�8Ϛ{!X��_M��(��U�̥�ϋ��T��w�k���.��o�~q�1ʷ��7[��^�v.n	m��U;�C���A�s,):��w _[X�O����;��c_�m��2�	�.��].��J ���V,xq��Xr>����s��Y����W�Q#Ţ`#��H �v�D,hQ�S^[�=�BΚ�uY7ة��9�O�,J�Jq�G��h�(`��a>����3����u��]��O������^$�O�|3�\������8���?c9�?uvl:��8�rAN�̕�X$L�����7Iau}4�t�R�bY�nUU�ͫ�f[~�J��"|hI�..S�R$���,�w�ֽ)!�"�������}Q�u_ڽуF�i��bS��ѳa�¿N����8〈�c��F��SC��ok�a(�.��B<i�x��Ԕ�RG���R�JEj�m��N- ��01�d�$���f3����lT�`��w��5F~]~�*2i�ya��Y��YJyo�.n�E$"7���,�KJQ'ւ����p���f���5��`��#�Aȣ)\Re�Z��{�l�����>P��K���p1���0>6j%����eAxkx%�>x&��@F��� �u���8Q��n������I�!�)��fA'U"�Ld��r����e��҈����=X"�zgH�y���Uf'ctp��j,퇰��2V��*���!������P��������+����YZJ�>�JnoUQQr�;������8
2���Z.�|?��@�_̏ܬ�\�	]��{���$�*�P� ���z�JP67qѲ�'����q*Y�� ����<�5?�p�}R���VA[}o�2��� ��w�Y5��6��2�q<&���>}�=��u��ݚ�[�L�\�L3�L	����_�M�䄬��#+)7���"5/�d�=�H�<7�gh)���]�@C4�#����l�,��M�z�w/J:d�p:3��ώ(-�6�*׭t4^@�>01����L�\xPCB�s�*�&ף�Y!�N��M�^l��1���>ͅetaNҢZBεS�e�%������ �ɣ@��r�.A
~0�%��Y���%<��:�1�bp3pih��X���Ri�%x�S�֨C�C-$y�eA^M��#N�%���L�Ϡ���{�Yk���t_g��ae1<�|j��[	9��b�m���ؒdV�hQZs� ���&"}15�.�N��́0���)��f������⛞��"��1$���QB�`55��vw��a��n��ֲ�{$G�e��������lr�.� ���@|C8c�~t�Ή�:j�:��L<:��d�EVЧRH�5%2M���wtӭ씨�i�Z���c��ΨM��Q���v R��"�=��&��e��~�L9E����$���:=�쾓͢j�vN�Z�X3$�N9�U;A����\�'�]T4e5f[��)z�o1H��;${z��o�a� �Ԟ��S��F'����:��󊑢�6�w��kSke%���̰AtԈ�(���L�#��Ȥf(b����e�ql(��KוdĒ�x��� ���X[!aĪ1?����Z��|� �����q���N�ف�.;�@���8������A;:�8���ĉ.,����d�Em_����y�RS�ssE^<����vM;2����[���O"1�@��;�`8��3�g$��sT���������{Ќ�o-iS��E,��72瀴A�ASv�v�}�Wm
����\�X�R��k��K �W:#٦����P���>պ-�};�=�yԑQs�òД��7��C��P0�;�ݺ�D��7
���?ūJGT+@M1�o6�<o�!�=TCE{K�������]>o>˲t-5�p�CįXi��d_;Qo���	�NZ�R���������5(�X�-��\���p)��y��V�e�n�p �Е�=�K~C���������Y5C�m2+��TK�Cv�z���$��V��e�vM4��e�͵h���Xxc9&P�Y�y_i~*�f}��M�v��	��AX�̣��EY���*�v������
t�.$�!L
�^:lG�'��c�dr.�$`�t���=o�z�l;⚽��c!w.�U��v���?��~��\hВ�5��*�2��I�#��29��S�vi��ł9xx;��V>ۄJP�[���_;��X�h�O�&.��ki��)�7F*��n���Z�>��"�(K�^.B\ �;��O�gu��#.���� |���V�����:������1�:B�������-s�h�EByT�շ�iZ�՞�k�
��g�(�vkn�^>>`��|���J�r)[}"�������������t��C��,�w�	�m��~��Kd�\ߛ�ĆY�za�T�����R ��$�ũ��L3
���G�����mҔ��y��iV���6e�8y��qИ˱�L�����\��園��5�}̫ј��9T7ɑ�/���_׶=�OA�HK�\��jN�R�#��G��ѯ�� C{�@f�������ZN� L� ��S��X��sr�=Pkp�נ>��e��ۥ 6$�p\��C�7�$�J�QHc� �4�!���IxS�r�^�h��@*,��C~>]w>0����/ ����;��3;��������7h��g�E���-�yYb���M���O�q�w��DV{>%?3�O�#u���5 7�.�1U|⩒0܇d��獦��PP�빺{�R�����_�VTk,�|�ob�y���G85��sA'���<�a/{Zfw���t��	L2�U�p����)%������<E�_�\���e�_����)�;G:�����"�#��PjP�.�c�!(��o�� Su$KN#H.q� ��8�����{BW##���2\�IA���}�Wt[]U�3����x�$�;�2(�Ƥ�-�ϵδ�{w��[|ޕ"]�5�u��yUV�29��s�l��L+(.A�p@��]4e'?�&�5�SE��&L��>J��n��t��$Ƕ�X"��)P|v�\7�d���ښ�fR����
��Oc�pr�>�0؂�.�.����a����pK� , S��Geף}�Qވ��	�0��p!�P`�������B�î$��
j�ݿu�aʞv���zl�:��z��5`���k��D�8O�U�U��c˴�X��)p���P��D��O�5�"�\��\9B�:�������K\^s�Xi�5G k�Y�snf���D�rP�V�Z=
��%ĳ��5Th�����Pt�.1pdt5�%���� �S�L�;g�1Yc�����<:���ŷb���D�FEu�\�CՊ��(�p?�^5,����Ihf�D��:�.>�@�$T^�� �O�U�̓ԻZpuO)�J�1����(,�M��}*��(�7��[N�U4姝�+�1w����#�����|L��w������Ou�!@4(�Ľ:��~�t�F�voXK��$#p�������J�
u��ar�C>݅s ~�����ә��񔶓��]Q{djA���a�j��V~���o_���U�B󵔑�Sě��Q��5~Ȳ��=N�[t���/h--��jQw��-FT>��?�Aiu9^�_��g,�E��)˵k��N^	�*J%X����Ϸߴ����+�P.���(��d�}up����?�0� ������a!��P{��'ٽ,�з⪈f��\[���rGv��#�ۯ R�@�e�>��C�Hg�K���r+����E&��&2$�t:����c���x��Id�]�X툉��lO���1�S��G��� �*�0��6����C�	�W�ș����c�������L}�ɸ]�Ag�V��W<
���<���
t���/ka�T^�5MBl�Tf)�}M�5�V�
��ռN�1�P�ל\#:C�ҵ�y���'|�+j�;�ؽC�րCs������v��̛LV%/�
���ۃ�����Q1��Q���;�%�� z����x�%�5K�+��H�g�#���Y�n���]�:E����L���P�2-�%B���)-%�e��2��x��x��AU��'�������{��`�{ϣ�}�V$R�����IĤ�έ��\�$�f���W~U��rs���ӷb佲�v����;�BH<^+I��3�tX�����v���Jns�>Ob�+y��&���\3�ק�Ew�ɡ]ȳUذ����xgF��~�ް��#��W��=�$�#������l0tT�>�=�`��(�G{�a����Q�X���n��8����M��C=V�m�ȷ�{����S�*l��ЮR��	%��sz���@��0�H��B�r��h�0@c��
���2n���Q)�K<7����O���j?z��G`�%(��1�wL�"Z	�z�s��������
u|	� �\p?X<��m#wL6,O�=��:D���q�J�\^��8sq3J�Td�j͵[�<v����',�g ���+��?���k2��?Io��|W�M��Ielx���r~� ��FWZu������+���b�q�Q:�4#$fMU�sR^��NL�;Ȁ_�� d/?d ������|��dv��z!�����K"�#.���\}u�X-�����re�RB!}�2"�'��SE.�s_���3@B<(��9k��1�?v�?���g�͜���{�bc�S��}g����?=z8[R�py� ��ᄇ�tD�^r��(�RTs�ӆ��mCm��:���
�$�6t��LQ�t2�'�����ʧ&�aa�[�A %������	���	Q2���Eh����̔<�I���A�q�=�Ӫ
�ba,҉'�	xen9��決��I������!�*t�o��4SW��jtC4��kƹ�p(����~h�D�nM��&b�\^������#8|;(j�ݗUu�R�;�1ι�nm"�?@#v���r��~�>�s�<��Œڰ�Y)�tz�|}�����Д8�}Ě�8�t�/V�&��D��&�)2��	���Z��c$*���d̠X*@
 u��gp�P�/n�09E�M��x��1ktط6�6���n���Rsl�z��^|��?�}4��9�U�L���Fa���;	ٽj��)�����)�~/SM� �n%7L�#^:Pl�f.��)�X������[D!�q��l��t�
����yf��g�',q�u>h*2�/��K��	I��ֲ?P��q�Z˱u����f�ɏ6	@9�p�y�Y�q\1��E�r�,���]�TBΙ�B<�b}�ޞc�f��Ϙ�Zͫ<�N�R�p��:�Ĕ84AQt�R��fXh�s����m��M���/w)T�͎���.�H��{	R�`�;�z�BK���O4T�o8,��n�.�q�d��V^4�Hx�c�#qd���E٨mE�\F�%�v�,�#S)ЇO�{T,�����xH����KQ:�%�c�0,-�b`�SZ�/�IV��w8&�ejC��#��/�\�u��)�e�@�o��W[�`�	T�.�~B��B��յjoj��?��n�8ڥ��3O>�{Zb��������~/@�(.�g��!b�e�H����=�2�����EA|�T���H0uS[�p��k�Ѱ+���#�/-�In�_�Ts�M���V�덷���C��;~n��׷�Ck���Z��sTi�°�b����Y�V�U�P8���At�kB�-I \RA�+=��5�� ����)3�bO2�>��͓__��T�'���6,�;c"���Cb�pZ~�,��v��3CO0v5��.Zf֗eT�	(�2[�@����H��D���G)�YbE�@��g� bb�&bC�j���Ե�3�J���.T�K���J�z��!��w��ҙ� Ѯ��Lewܛ��jɲ:"1� �p������?�ci�-v��X�����;�Z������J�~/J��I�a>,�X5q���}s��/�mq�:�u�y���`�oޔ0����F��oooEA�j��m��T�ې͊?ˀ�fo/��KN!I�[ �j�q�1�^7e�k�٧����0�������
��oH%��)J��e�}��x-���k}�
>��YAвV��#٣�B�6��th��<�<R�~���3�!�H��H��� ����fP��n(_�����<1�)���,��� qx��ru����Z(���M�²2�썐&��\J]8a�9̩,��I%G��@,��H?b��W#u�9�S��)[�"V�x\���}�ǌ�in�#[R��[�xq��3��DX���f��2`���P�e��rq8��1ۼ���A�:M�#��<,xI�fz�F�=�,����x�����ʲ$H��؊J����kQ�M"rf����W���e�V>�B����7��>	��tU��'610�-ŤS���l�ĭ1����8�}=fo����3ʎ�3�(y�Q�?N�C{�<eMh�#���)��s�pP�kG1y�me�B�l�\<�2���iS���l7��W��fA����:��ӥV���N �KJPk�?Jb�/�k�e�(�S:<'�(��۱��ϒHH 0���/�����3i��6]�m��@��#��t>��|e�q�`'hZ�E{8�{���M��@�7$K8pF���L�ǘ�Tȶ'�/V�ޤ�-`(iȕ��-L����4�oY���e�>������1�zx�yN��R����JL���!�Q0uJ�����"��rKCj@[	̀���Bݭo��Ϝ�߀�L�rq�	����k�^�>6���X�鋉���|�Һ���H�fE�Sd����2_Zu�ȧ�ӣu&b�r��#j�Tկkq�s�?ָ���d����+]���~g�s�?m�(+t&�Z!	tvܜ"o�1������d�o�Y$A=��.]#���V0�<]��s��%:���&����_�pI������R�p����8��-����=��	�ه;A��w���E��~���Ψ����`�A�`]|����Lo�yA�!CI�dsĥ�}���V���ֆ&b4 ��}�t[��m*Q'6)yh� N)��m?D��ip{�ѥ�/w���֊�ܜ�^��CZb1�u"��9x/'X�B�������=�-�|o�>$Nf��{B�/�3�Ěz��+�x�]
�y�:�{��l֙�^�A?#�!��y�l��p��ؾ�Sp�=�����{�bH�)oBnI��r-e��=<���gV]d���<fĥ�H���U���F�8k|��2�/���f�Xe1�.DEIǬΓ\��ŷݔC���d|����k�N(����Q+����Q�u���8<5�I�~�m������f�� ��C���gsB�* L�2k	�X�8C�^��g���-�v1,\p6=�Z%���[?>V%�������z�>Ѵ��B�~+��B%M�`&ow���w,lʼ:iKJ�#���}WL�Bڨ>��j+k��YV^΄�I�2�/�݅����p���0|;�6��G�Q�N�W©�r��~V�F-OCK�nw:�!	�kZ}_�AT���I!�*Ъ�ue�-�Yw�6{:f�-��o�G�,����~G�V�,)�GP �!v��'w���bf�}9wm�l�?h6Վ!,�Nq������d�i��Њ>/���������i�m�N��j0�(<����Cw�Y����0�iik�CmV�}�O�m�X� l�QP�CR�,tW[�)�'t�h��5!���=a�\�C�Y���
8I\��z&a=��q��̍n�,��T#�`1EZ%��߮�;���R�ᅼJ��'n�]��Sj�GK����?^�o�Y��9�!�������`��	�ٍ�SL��P��`�AY.��@xz�����5�G�.��6X@U7�?��vU�`F�:!8_@o�a>��Q��L��u�X�Xߢ<�#��~�����DI�F�C2���u���UO�>gl�;K�TP�Yw_�n]}�L���٢����S"��\�@��M�".H�/=��bc����#/���H��
��/,��R����J�z̮�=Fa@qZ-��`�����!�yW�dA��%Yg�Z��=��s{�b7OR�ÛJɒ��uw�O���<�$A��4���Z��68z0c�?��!x=,~2񔏆q�}����E
=O;%I�m�Bڱ�Jb��tA�mFlU�vh�
͓u����I�Ϣ� ,lVSnp?i��[	T���?������J�^/��]r�.8�BP�Z�.��@3��4�� ����Rd|X֩��"+n��XId���#�P)[�у�4����;��au�41�kG>�`xA����_��,�ND��@%�I:6��P���y�"s���p��<�d!����i9*N7�B=CA����K�i�����-Bō���;� �$��Åŗ��M�7��(����V�`9i�a����~߆���������SvK�@�(}�)Lxtg8P���6$���>�n0X�Y�H�~P��?�����IR��4q�x�r�@�lK���s�{Pl�n��� H"�$w��ؖ]�Lz����,���o7�|�?Y��c:�'h�ݷ��%� PI@ �|�l��$/���%�P�	ptQ����(�޶�i�+��l��Q���}����I�=��E2ߞ��P�|� �D���;)����YP�\D�ɹ�Hk�o�Vww ���P��0��}��f��X<�(�@;�$������	:��I����..�?Hm� `׬��wi�^��*��>f`�lc]#�U�C��z�LJ�Dion��	�,��\�W� �|�4֋Ϻ�q����i)E��W͡���Sj��F�b�"�Ī#�Xx8�.�(��[ ��{o,���DЯu.c�0�������T|%�kM\��Oi�� ��rf`ʲԉ�c���g	N}�����|�˩���v�G�w���01h�@S�q�;π_�̧p?��/7���,��E��F�.�J�s��?�-�Q�X'��7<���?�_���J��*Z�/��>�E���ʸ�=�g��/m��4���z(�@�[��f�E�H��L��)z�����s��{_��Q�1�w��B��/�	B�6�5������4&�I�9 ����ς�������iO���@_!Vw,Y+�����{<T:?������?���19|�"������7�>�����ѬĂ��7 �Wg&���Z�����xf�P5�(�ݚ	h�����g��vO�3��.t���=�
���zW?��m	�"R��8�fEat��9�n��spuw�t�r]��z�<tM�"4�_*���W8O�u]'߰��d>Ғ6؟�<b)�S"�w�ˆtpI:ܗ2���")Z�ZJN
� �,c��#Orw�z�q�0�~�餅e�AI��P%(g&.��o��]'`�^�(P��+kZp��F���f+
"�}t1Y�{e�4�,�*��݊Z��:�x׉ȒR�Ɵ��<|R��I��(������>m���LEa�$�?q��D��W��1t�M�~��/�.���Ij�B��F��X��}R�.�+��G*ևIh�xD�OCU�\�k�M�XQ'�=�J֒͏]y���5�w)���#�����Η�y�P,���Y?@�/ĤN�q�XN�_Qh#Aw�"m�ؓR��g�Yַ
粚0�����ń�/i��O1���[փ�7u`G�����?�o�U�rYUl�>9~��x'ۚ��)'���d9f�l2H������"���M�)��̓g7��.��5�'��"k��&��>\���1jBe�!�,`N��i����><8��tL�����&4���[^2�f����Aj���1����<X��б9n��t��T5�2u;��%kKzz(�fs�Z�3������H������C�fJ��pʆ�Q��*�De�Ǧ�-��Q�p�^��V:Z���PY�}�<����D��)�'H���g�������Ç��eB�mX���D=�N�M�s��|��-�M��͜�U���TIKc|�
ŉWs�F�����?b�D�;
�6$�����$�fogq���~=�Θ"r�VTF���4�J|����C~��l�o�/����)�}a�Ǎ.4�]���32N[�c��Ė�w��sS玿;5������2O���eU�����V���	#L8��EV`���.������V%��1=*���=8_���Im]�� \-i�N����X$$K�}�n���ZRB�$'�M5���ӫh����ӥ�EY6�hx���;�{�[;���wx�e�8�ք(ԭ�g�y�u�	�J���th�3��O��Z��_	}��8쇻�!�/Qj��@���}�Q���4�0�{�sc����q��9�����R�WI��(��Ѷ��9��`
u�KG	sm{�b���񨢏�}�T�y�!�IE��/�	w%ͩ��{Le$�[��#R���a�B��`�r�Bn:I��|�J��䴷�RI}�~�a*��/�I2��|��OwO��@%!�Yf�"8�b�&N5�u���o������r����i+��W�����e�Z���Jv��8RW%�Z����͔�8��'�V ���;��I��L�-d��\K���_���k�ӥ]��{��#���j����c'����l��s!��%�Q�������$Ј��0>`ʖA��%\�[����� �A��)��d��"�]�(�IRc�#f��nxy���h�R|��7;�7ՙ��O9���C{�����)��ԘWS����[��4�>b&�j��1<�_��x�.�e�"��R{��U��&y�5Y�]FQ[�Z(lwǡ(VH�7�d��0@�^��'D��40h����̔�v����M��)��rB�9��*U�+�Y���HAԘ,Z)�S�D#ؾ�ľ�ο2^��/�x��`� � �A7�.�;�@���&}� �:�	���&@�\x.�L
Khr A���FF�o`��@�8����D:�����f6F���޶Rfրfy��SE��n�;�IKĉ2ؐ�bUlH��"�	n@�;%��'�&YF���4���YfQ>�.�=�송X��Wk��0o�f�T�[��[������b�;8�m�G�Pb;q�ݯ��G�/��؋`Q���b�q�̖{&8 �}����MOxG��m��a��4>����
�'�lL��Sj�#��_~���;/�n�ף�2&�5�:���$@��O���jqnM��7�em��v
`�����RCu�|vI��̲�9��5.!��7_�h���I�xņ>sra�
R"}Ʌz�-c���p�<�cp4��v��å�6�����Cx](�7��]R��j4/z\�	)��6��u`~��-��\T�q��H�#�y$����Gk�n��?�/{��w�E����B���:���������4#!8l
f�+ �՞������+���K�	��'ͧ���Iɑ�A�g'}��&��\XԆ3Ӣtҹ�\n�i�V�L.!�i�����~��N���RKv�ׁ�{� ��iyݮj�^��va��)a H77ɱ7uC����[ox��w�3rז��*����F��ư�9[ıee��=�������Wx���?�w)gݣs$��μ����&S���\�1|����>F�\�a�7��#f��B�[t���Q�����n1�������6�g�{z�>�i︅ ��Ѩ ɦA�]M��r�!K������?���/���0ԣ��E�>6R#9�����Aϵ�P�R���s��ʂ�H�?<I�nOO�`�nEDE�!S�@�K��͓��?3��oA��,4���-�Ğk��z�������=�G�ԕ'g��Ut&2Ŕ�KQ���D�P[�*����G|	 ���&����/�n��o��}i:jc`�_d���9��!8�^�zR�	�	d�Q��܃f�] ������\n&o�g���ʙZ1IYv���n��L��)
��v��y��?�켑�	����-A�0�|=%)$A��E��}����z�W7f�K�X��"��gw��/>����O�$�G�C���2O��M��f�l��dN�DD�1���Uk%3�o���g���m���N��0��� �S�H*�kxShi�L= �o����mME���^�������A�↩�RM/�s�������ӈSLz��)# �u��z���okG�3n�QB빇Gp\�3Ɲ��x�o��@:��RT{Խ@�Zb����ԨDP�W��f���;�\��l�Hy92ہg+�=A�T,e�:W�?�%A�ʌ���y�نsB�~�63&�8�*M�En�O��+TYf���襚�o���HF��U��5�j�� �B��n���LS@�xP�Y %SA�8�d͠g(�u3�٘^F������E��FA��k��;a7
:8!�:`U�&��j����u���z��ܣ�25HR��ז�j2�[F�|�v��/�8���� �E����~5j�����Ut�R�rA�3o��RĽt`W��e\=� {)���+�X6�y�^�ڛ��[3.�4$�����S74Yڂ�{������F˘ʃL�AF�_�)l��&���L0�%�U�1_@�<X��M$VN`��]ܙ��}�sJ�e?T�st�gg�����7X��|; (�`C�¡>\UK�Ŗ,S�~�c㣔�$7'w¯S`��.��«���Z��ċ&L�3#W�j[�K��k��Aʲ��ֵ��`7M�>Z#K"Љ0�P��ҥS4w&F1r�rz�G��^gn#�}#Ժ.����t�ʴ}�LՎ*h���F���zF�? �i̦����(}�	�}!��k�� _2�U��I8�\֋l���<oz� �}�"����Cj��.�a^"��"0*ݥ����'��	ay�/4IM`�K-2�Ͽ���#���Pi��v�Q�[��7���w�9/˱�aj�N^�+��HQ�?��ڐf��V$���-eط��x��LOB��G��:4� ��Gm�Z��ywvz�+�}�$"ecS�	��� �b<�XOvO?���g��U�v6�Ċ*g4C��v�D��ڼs�	��7�+��x�I����G���3�`��<��;���m�#a�.��d-c���A�b��������][���h�7��pf���Ǆ*���G/ήuX��\��o��cr���/�^���
�0n���7t[�[��<p���:�s��H�ᚣ�MXe�~�l�;d���0-CC�|��U	%��:�K�w�"�x�gWDsG��u?
3��v��KķT��g���陼�84ËK��Txem��H윎l+������E'B������j�wJ~�す�J��B'?i�)��Em�fߎ? c�e,G ����� zr��l�F;����6Hۿ����L��\��,��}�ۼ�&<�<�-���JB�� !eL(���"�K;��v0�V.RІz���䅯���ڇ�Lc�n鲞�/W���~ H��T�����Z3}��g�V`�ӷxz�Ab?�4��Y�����|kA��6a�ܡ�q�_@��3��ŝ��
0�T�y��"V��uZI:;����_l|�)��W�c3A��f�C��k�ʿu^���yp�*gBm>�!XI�q9�Y�������W8� ��4������i{n#_ �դk�6�,���?;a'���?�> #�K��z���>����1���*��xo.&c��VlYy㯭�_gl-(�xd���=~§��
E�d��8N����3��)dƮ���i��6U�|�[���La�`t��QTQ�:��� �^�� ��Z�ˎ��E���՟Q��O���i����l���ۂ�Ԍ72�%;W����Q���o��~�"~�:\Mr���a�7�2�"�9.�p�	{qQ>�	q8�E͟�;n�O/�����v8YG�M��Qt�@�Z#��D�nA��j�[k�С����Y�y�V�Z�ҳL�/���	��d0��/v�`�DR�?G���'ޟ*�Q�;Ur��� ��'׆L�
�.��eS$P�.��X]q'��D*H�&@����ax���D���ѣ`cj���$�,ڗ5e�4�נ���c����a���åj�e2�Wô��O��׌��u���3�nd���R3�i"���_J|�Rޑ��ZN���`󜬀�iJ�&��\<z/�Y$x-���j��f�t��r�$���`˰��pFo;�j����eE�'fCW&VU�h�������l���t�[SE�4~�\T�r��"��A��aET��YO�Pr�o�Z�̓u�����?8��uzMBN�/&� �� 7����k��
~�>��Yڜ�hV���r[���:_msJN� qN�����P�=�!������=d}��=~^|��뷏��D�H�Ҟ)?��s٨h�#�ݪ�׷'a����N�!�������d��6W�J�c�W��E5Ю?�<�> �ˋ��(���|��$U ��qxY�z��]M�.f�<� ��Ȇ��v�,Q<Y�D�Q�/�TJ�Y�t��jӏ�V�u��}�`b�X�V{ T�HZ0SUYo�0X6�oe��	�����\�Μb�T��%����y��Y������X��g��j^�H}ҼS�ʉ�n�1����	��d8��$k7�}e1ч��!:���`�cy@�ݥ�<S�iᦞYp�8/V�(5��R����Πlh[���w8;�M��]"���6Ȍ�����]@x:̈�/��B4K�
zTP�o�����ܺ:R��Ac�ĭy�����1�]�Όv*��X�v�O��d���vjF�
KJ�x�KR�K������ɐ�6��������PR���Ӊ�����lN�l�eL���L��:����w��c<,s1)9�����=I���u�uwv�ו��o�T}稳�����1�ݢ���?��R `�xLU�V&��?�曾K.�Dʵ�r�	����H�Ś@i�#Q[��Y�B�ET+�$'92'�ͻ��s�K�Mm�����a��o��ˎ��"�z�����$��3�Q򋡀��ά�s�9�lތӪ�76��%�eQo���<`1^�D���jR�2w�,ckW��X��=1 S�I�J��j��,aϡJ�<��WZ��j�T�ޱJ�UL1�) �0�?�å�������-��I���b�K���fU�MR���p��/��J<d3pe�t���1=ԃ��ĞĨ�B��
�6
�&��/z�st��x��k�H�g�O���U���l԰�� w���!I��e#�u���;9�����(�Կ�x<�#!�x[Cخh��mH��*U#�3��t4�A@n#]��Lq.[V[Fu�i��R�	Th��DY䐧EG�'E��7��J��CltN�5`n���cU����1�k�:)`�'�z�r����W��Gz��%ay*�p�	-���W@g˫�a���Gm����nX�1u֑d�f4��4���Vᨤ��6�g�ø��$��/Ca��"�?ԉ:gĞ#3v����2E�,)/����*3��Uc��=L]�#�sѫT^!�"y���FY�d	��;H����i�-�pi�B�΃��3�%Sc��]@(m���z���Z���ݯd�(5�p(	��mt몊�y�����d��wN���G�G��ƅe8U�7�w�:�:!w�=і,3L�v���{m�������k�<�n��0"Y��ǚ�u	|�P�_*�����-����r�t�Ih�K�Ե��*2ƣ".�(G��i��ɓ�T`G�2���&��N����
>0
#
��]=�)�~ڿ�@�S�Anю���H�����Q�sԻ`s��b}����a7(]Sk0�~��=*#j5jj!�g���i�2a�W�=��Z�|�	�r˚�N��X��Ǝa%+&�����2��^}��$���j'�h�
[G��J�|#�[�H�ok�:���mݩ¸�i�zN�P"D��Fs���,��+ӆ�)-_Pt���n�B�b1���G͉��,|�K)�	V��x�*1�y���V�u�������?&	�w�5f��kc�4�]d�V��}��l�<��6p�D��z9��C��� �&_�H�`�;����x�	���gz0y�~��?���ChE���ߡ�k48u�T;���KgJ�i�6�v���:�Z�^0J"^J��t�SpL��o����iVg������ߢd�]�8Vk�/,/�Ih�犓B��Y!-��0��!�É����#��?��{`�
�}EY����Y���Y]>��~z~��ȣ��Q���Wk�F��`�N�k�j��oZ�M`X	��v-p�xS� ��8<V&���卆\tk_P[a��-���+��r��`�K\?}�n|c+�p��)�o�P�w��?���id��w"�(����,u&�B�b?��A�}]zb9��H��3����v�g���_����9����� �0c�9c!5����L��j�Z+;<�ٶJ��"�`*�'>IO�oq������s�(mW1��1��a���֓���x�AH�����`'A��^1��q���W٢�Á��.(8&�[�xer�ٌT���������&��e̤0���w:H��e(`͹�(zr�|� �;-N8��XЯ���U�a.k�s�����O,���
S=Q�g�D ����:Rߥ��w�ٝ���2bE�נ~W��b�a5ŀ=��������N	h����w4t�V��Z;�1_M��Xo [}�v=�o<���u�	�����ak2�2!���J\&u��wAڛ��δb<``�*�"A���3u-��C�綆��W��'2�
��@_��^c\3O���Wp��aBMT�(D�x��ۚ�G�9V��(e�P�����K�&�"�v4G��0|�\�{�;X���S��5^}�:W���d�j�̆����r�_��8������o!1@��+�í��i�����?J�ը��hD�"գ�h��uW����"n�NvaL���O��Z�}.cm�� '��16�tk���)��u����'�b�d������޷�5����}��c3�/���[)� �O'���uh�{�6�\O����O#Y"�r�e����.� ��@���s�Vr���{�{S�M��t�d����&#�~����!������
���p��%Z�n�:=���J�f~���c[�������$r�����H2�q��A��I����5[9R���/�S�&N1���u����/�mͦ�~j{�#������{D�1v6M�9B+HKNI*1W��z���hkƌ�2�*��e���dpI$!�D����|O���N#��҂jY�c��r�`�~�b��kP/Hʙ]6~�`E0���X��[�^���$���R?�J�i�F�d�xh�)��5zc̕OB3�*�W�YS��7p�[�Dqm_�x -�_��s�s��k�����P�l&�y
��M���#��b�|j�V?�x��P`*ƣ $�/K��ř���n������U��$rA��p�v��./��S?�mr�In;����A1Etj$-/I��;�s�/��35'�����O�C�:�����Y��ÿ�]*T�\�h�=��#�I9鿊��񌧛k1�=�NW�)q�U����ē�'O�%�0��a�MTaE�a*���__e���Kh�һ.��zYw�ʠ$%��(�Q.)�(;"(Y����h�&=��"a3�@����JCryd�*f�(-!*�mx�;�����r����e������t�ȇ���}���{�"E<���$�s�yջ���I�=���(J@�,a0�-Ǿ�l�F�W#�ϕ�((��0�����7���,�s��Ԃa���"�����@MEcf��[���G� ��yPx�T&�V�r���������!OM���\�rZ\3�5F��s����E�!�[��"E*o�ۦ�u<��}�������4�R3����2ۉT�������uPIߘ�p�������d/	F�_��g]�~�?^]%7�7�Y\�q��(�^�喲@L'�=c4F-v,7:J^��t�B����y�}e�����mJ���������h��2��y"�Rҝ!3Bk�K��G���sz?LY��	�v��D+�����z?����P���G�G�|@�м΂��=F�K�om�U��0\�����?���^RZ�y��Q�,��~�e�\x��!�^�X�IjW�u�w�4X?�c�i��ra�$�
���Tn�5f���Ic"��Ko�0i��J��w���!��v_���������x�I�_LS2x����ϗ�Y�=+��
^��878�;�x7�ދ:�8FQ�A3�����b�z�@N����WDVa������?��Ǭ��jf�օ�a�f�m�_��p(��<B����^&�!��=��9��:<�����-�`s
���"�s3�%�1�2�}v<
`#� &��9?��!1;��5p�%��~b�k�ĚI��}��h/L F�8��o��j1E��I��Ǡ�F�L?a)�>�4-T���O��u�ҏ��^��d:mc#b��uJgߒO
Qe���z����wr��i��q��s��=s*c���D{6/����)�8�*r�ͺ�kX;����`�����@���RN1��l�w�Pa�M���<��X������#�?G�S?�Z�����]���\P3��2�8���/G1�>�F_�ho�Zի�y�*�����뿥B�o��N w��4�=�� ���¹�2���_���N�f&$��TU�QL���2�E0����`:�uV�Y��+������\�	i�]B�:;!��J��eN�}�C�;���fhE<w�;6;e���'�?M����vc�*���9��wec��y0��y��M/%�Qj�X�_�,r����N��l8�:�r�Q)TQ�A'�`���>�'����0�g��;)�R� ��
�_ ��_�9���"�����H"/��x儢_�u�2E����=\Q�m_ # {�X��X���y�:��!�Z���G2�.�%�/��;�p�c�~%>��(j��������y��UcBr�D���h#b!�Z߹��\��ίh?��o<K*I緢�^�t��IuLX=S��)j\�"+R�A� ����&�﫷��6��t��)x��5���ïg��d�>ݴ�� ��>��V�S�u�pg"�`���K�`���ߛ��Ώ���ט\�^)��V5@�Y� :0v��ҏB�5���� �*�]$&�`]���:��&��_D�a[��EW�������6ɨ����C�3�=�I�ѥ�|��%x�c��^��C��l�ʏ���~�z��~���-�w�25p4�DBw7�u���v�����,4�=AfıO#X���pk��A�$��1�f��z��c�ؘg�������(����q�)�`s�2"�!��i�8�^�n^=��S1�j��i{Nβ���~g�fY�۔T�[Ж� ]�w�������n�\�NIIw�$�n��o��}�1�%Ae�*%Ѥk�=qC|�Z	�6@�غ��+Wؠ�)A��IJ�D��4���(3�ȆdQ��{xƂ(��j�X/K:-��=���},1u��z�z���v�|>�ү0��F6��cO����h\���.>y��P��OqX���8���p�-\,U#d2+w�9�=Q#hQ������q{���)��L�w�N�i�MC�<r'`@����,{�1g�ΧIl�C��t�*�j=�H.�}5��{��<�"����F�u����`w��Һ��ıtuZf)�$�v�a騦�7�y�Ee���������_Mh[7�3��IC��T��]�V�pt�zW&o1C�Tʶ���?��n8s�4�X���p T�����Kͼ�����G�@����[@�5S�qJ�[��AR�Mr���6���Nc_ȸG��̤�QhZ^^����k�|��C���P�N�\�m�o]��K�d)��)���ͬ*9��r*��ӛ�h$Y 3*տ*yn}���0o��[ey���hG<�ҙj�7�L��
 @v�d��k'C"�&�%ȿ��QK��-�����ଂf��qQ�ո�xņxν�gr9w5��ı����*�n���r��'��v�t��D΄֮y֙������D�n�t#��{SPhB��k��2��j5hw�<C-�|�e�S����t��v�]hg����4.�C��)Q��XN�`_eq�@��U�P����2ժ'�ą��L�0�_���uX���'�:��&`�`t�<��<�B�u��Ʌ����WNO�[�AH��]*�����zCDcƣ�QKE f0_˞f�(�;�?I��J�	p���qa���-�?�u2��̬PX�Qg��s>d���˽�u��(Ʌ�n8/X�x�2�H ��(��Y�@�:�����ZQ,��#�ܝz�	+Q���n?}�c����/-�@���*�I�-vMH�z:�L�w���$a��k��?Y��cS+���F~`q@!��Gp_�
�ꦊ)@�cѼ���W����]�w�^*;J����E��;j�R��$�������Eh�����xm^�h_5z
���exC�Kr��hQ���+�aZ �±B�W9��E�x�b�fPr�p�I����[��aT�uM��ڗt���|h@��!�NʞW>[�5�j`��vo%R�V.�0�4_���~�/@����)�ϣ�)��@�malP���=�1�hQ6��-���Nz_6?X5r]�Zyĩ+��]ƊXb�v~�p�쬿�ljY	N��Tjՙ-b���χ&XG��;w�8�ʞr�H�%)̯��r:�D3�A&�Ʉ������E�Y�fh�z�`�!A�m.�;]͂�pr�Ueݟ� �p���Ln�������^�����9�)���b�B�P'��
>�b�&Va�Ȥ@I�w��-8XTi(+*��ILx�I>�N�l���=4z}@�X����w`D`�W�Q�J�2Y2�w��Q�A�H3S���l��RF*��FJ���9˽o�s�vKVJ�]?�zCh}���!�+�*b?_�.�3V�!�w#�_��|%�W��>�Iw~�KY���������.�=1^��Y��i3@1�90����M �>�:ɔL�0Q��������Z�-N�/7JjgM��F��<��ĉ<���\C� �V���k��ц��1Qӌ��у���'5(�W
�}�n�����#�T�&���DGsHCp���<w�-����P��c��*�#�?'�����@
�s��tB�R/}�^����*,�4�(�@H,�}�j���OѰ���ź�^$���(&:ۅ���ɗ���H��NofOA�j-��ps�$n a�eqNcJ�ü�V©]�i+I�Yu�eǾ���L�X,>Tr�V@_�
����SH��x�Z���'�C�EMY�D�����)���`E{��]Z�/l�q��3U{��Q!'�����u�tA��j=Z��#2u:��A_��@(�:1C���@.��{n T�KHfZ���r#�T�Ks��;�
�lL���H�bW	%$\���y�!��W+ޑ�v�M �]Y����
?.��f8���ݻ9�<��pہ"U�ޱ��k%�O#ڏ������I����Eh`�s����p�X�&U?�m�/��Y��k�(�i�T����Ԧ\���e���qU�h�&<~�����ݕ��_P����s^��D$�]�	���H��wߥ�6i��m�i��xP���rK#�i�z�X8T���9�o9{�=��uSϢI��ލ�Cc쾰��DP;X*Jki�ԩY�Cl+�mmȉҫ�D��]5�����T~���N���hƼ����#$T��ދ����HZ�^����a�`����ǐ3j�àt������o�!�ME���x�ynmĊ� �dN��%E���	tJ�a�������d��)����~�n�C�J��H�ڇ:B�<��O̱�8�{� ���S��"Z�-郀�Z�c�����e�ڢY�rUm3〢�VitY�0Ԭ�$���Ohl��*��6�L��&��I����H�q`�OJ��G�N�L�˸[�ڴC���'=��؀�0ΰ��3�4m�0��I����ۂT~��,���?3��!�%�;2$�}ŠY-i�)V�����#�ix����q�:�z�O������D��b�;��w^���.c�j�@&%=;���M��6�����ǜbs[�A^_������}�p�Ӑ���r��,^C%}�k���v[]ݽl��"��72$�0���:�,u��
�;����.!�&�.rg|������G�l1(P�T���G�[7s�S��%h�x䬊��g��0}��Eq�(?ں�����加H�T��h�5���L���>P8�ss7�������ۨ���j� ���ץ����xh�SwQ�,a���S����H���Mĕ�Y�D�$آ��/����l�I��>�)^y� 0�ˎ����_?_��F��I	u��F�#����敊��4s����,IP%����Q���J�v�,&�=D5[����.�֥��۟��?�u���~'���E�O��.�|��^��f��Ϛ�˟P�� �3L|U;�,0$g��`���襁'��j��ٴ�i߲Z��OJ����b�����<6ch��e|�mGͰ%RUk�p��-'����v� ��;������C�E�F��P�������.%B#Ա���ȱ6�zư����>���9���U��\�����Cp��#�y�F����W�Qcn/� �����nSTŽp'���06D�D�\ �y8un|���Qiȷ{-!	TYe�f&�93Xǆ����${��	�B��RŒ���=�?w/Ph|�Ţfy�q }\���d�-��ҢkF��=��oR�-�c'�p6����P���9��^V<�f��[��I`(Q�t$�n�G�| ��P��PP_R�͓Jr�I�ɀ>Y�싑Jn�m����sfɾ���_�a��Kzm������j7�`mH�6%$]S��`��;#9;�y6�;(5���R�my�t8�X�)��k��_�:� ��R�׹�p��xS�������纝A������a��B�C�G�{:<�n+%(rS�������wk������|>\o:�� QitJ�q>��g�u&�r��I�";���a2����ƍ���P��ڑ��Q��|��}=�Y��'#ێ�饮;��;���yہw7[�J�F��V|�O��~L�
�p�D+�7^F��G�%L���)��kwͱW��n o�zW���l�f)��"ޘJ:��J������˳hէQ�m�q俐)�x�nw-����_z��ȳ��Y9�������_,xn�v/2J:�Ŷ��(a�>��heJ�����T�h���\)*WSi����z�7���t�Zqs����-Й>ӤʈJH��3�*�#�{�5��).i��)��jU�7+�y�g\+?�r�+�(e�bc�=R�B#_����e��j�X<қ'���,�l��Z��D���xW0��0�W��uD�)�u
�B�D��)6PEسC%Q�tu�932Sm��^�W�%�ԑd�����$Ot�O�ֲ��<���Fμ����f�2�K�k�K��1��	L������
���`�*�'�.��d��m*8�������֔3е<a���e�ba_���dV��@Qϓ�\,̯"�hZ����٨HE��!�����E��oI��Ŋ��EMʹ2mgle*����F8O)��j��V2\�s}���5G1J�}k�M&�D�
�g�P�'a�&���q�PY�Kf�eCtwWzOY<��L��P0��Ą�a����*[̽�S[�� ؙUb�K�n����
^^�i�L�j�t�Jg�������������l��nd��)�I��D�a;7hW�,�y�������Y=�����';����S��Bb?l���͙�4M
i���[5L%jG�R��~ae�����[��ON6M�tr���SG��A�5[Q�p��ޝ���-����{`3a�gh_���
^8}���h��'R�
L������t�j�iOQ��E��>�J�,KÎkU������E����rq�qܛ�A��ZX�ެȞ*���C�ξ&n��~�u��RrE����mI�(ʢ��h�.`�(��:�*^�wh��^�Sm�y���S�f��p:�٫���*�a-ȓ~{��i��h�mtp��3fП����vW/N�E�.�DY絇8�L���0�4ÛF,�$�Jm��NE��_��/d�z�nK��l�y��.���˅�d0̫�?��J_�`��i:�V.8�"^,h�ǅ�.)b���]�cȦq�X��4vN�1?bD�r��x���$aH>��ߥ!A�i���1R$����:%8�RK�~��I�KJ����+�Mj���D@>g�<��J��N�-eq6��6ٟ�FE�ӣ�)2(H��k��i���q�?s31��8O����u�x<��m�jߝq��.%4М=�{�8+G7��������  ��ZoIs�g���b�_^����'��NO���I�X ��s�2�>�P	@Ϯg�,:�I�2N��}��Z�w��6-�c#d��`n�x�����	�+Y��l��=��1$�v���Ǚ�*��'�{ �H�-X<P��3��{3� ���g����~���/�o|-��zK��t܊w�7F��Z� ;cei�W�7��?�]���C��%i��*"�3�@��vo�{6Xe��n�F0l�ϼ&:vA��?q����38|֗�!���8|��һ�Cd���Ν�Cp��\"��2�8���I�Y�"����(�?��]uK�B-\Ȉo�����wIY���OʳD��7���>,B���=a�5������+2כ�!���K���*P(ӕ�v@c L]M{�:�F'S*�{�^L���W�{;gFb^u�p��ƫ�{y���4ou����~�-/	̘̕�b�_Kɟ Fy�J�ϑ��ρbɾ�r]��;�j��IoAQh��3zƒ�m�%�aU���`�񳇘A�4S3��,��}"������5�?}Y8V���\#_>��S���сE�L/�g�����u��I��#�=X���Z��jY�*V�^$��3\�g�Y�{�6����U(2��,�w��աޒ[=��1h�3O�?L�,C���~i�� �2���W�\�`��3�%�~�R�B�|
M�XT�5�m���k�a�4��|��j3p��/����"D�<N��p9��C �;KL���-��&��[M��2}�0o·*�:� �M�5�kq^Ʊ9C�#�+:�1^�8B�sV���cC)����n�����ڬ������������7��m%�ޱRTDwlw6�O;t���y��!* �=��c�G
+2�Z�'��3�˝�n�Nk4>�6KI��ïR�q&�c��8�1T.ѹi��kH�E�a۩9d����7��dK��7���m8w*)y���2�[D�}�� kFh�\�f����H�ϝ�9b���p�,��:��Gvʏ���18����1q�Z�9�8z���i/pg�r�+���Or�^F6
#a(
���cܦKV�qK:`���ƛ�s!׷��q-Y���ށ?��W�/�D�)n*B� o��-d�*���N�,��e{(�s�	�]'�\��:�wlW5��HZy��"�N\0�U�Q�7FȦ�Tѣ*�NO�TM�7��(zm4"��I��Z��웩����F�yq`�����x ��xuz�����tM2Ԥsu?x0�N����
���tŞ\��X�@|B;�D��lnkPNr�CjU��^���u���R��&�_8=����xebNɸ�YϽ�6�^��& �Eq�!n�m�;�W����|���B��:�FÓ,�* Bsx�H�[���#��(���y��BQ�aO���0�m�k����<�\쬷z�i��s�Ѡ3�݉eW<	y��n`:n6����g�p��$��0�� !�.Y���rb�~�i�%�����_��<��*�(��ۤf�L*�ԭ��&�۫>������ME�%����g�;8�lsVD�Z(D���]��(ax\������n���l>k�eV���6���6�\Z
�d�1i��e�VJZ4���ǫZPd�cM�fDs�������]��I��wn�q1�"}���\^�K5޳[Qng 4�]k����/�3�{	�"2�?���?l�⭰[���M.�<w��v!>T�E��{�l*��]71�^��w �����y� d�@�|�^��y�/���J�4�R/�O[V6Pˋ�a8������}M$ҳ`~b��kY7���j��x��y?rb�q�"s��-�=$LG8#:�P��1 _���!�惕b���܆}[�����`mN׳M���h��*��'�w�Ѩ���.L��l�&`���/���?�d�+�_��@��4�����q��_��4�ޭ�X��{�m���1���H��R6n�Sr`�zB\����l_�{aQ@�'-'�]o��ŜM4!�U6��n2�<�矺����Rރtgp+���ٙ�f��x�z;z�5;�n�'��m�3�l��c��|ސ��Ը���O�*���<���=�t���3r��j����K׊�2/*��rt�z�����8�P��M=���G1W���	YI���2N��
n�Џ��d����si������۩�2r��gQ*��%P��p$�Q�����(a=�Sx����A}�s3>!4NKHP�x1qy�$</QQ��y�C������<s�tT��fP1�ܷop��.������U�};㶒�R�"=er��(��1qO�����rtC���b�Q<:NN�y����^n��&=^]���a�jv����/j�J�0�����[�N��2��O�;�����cX�aݠtOh=��.w�7-�e�7�O�U�_���@�����8B/�z��Ӡ��Nu�m�܍�xF��^����E�H��̂(��@�.ePz�O��-�Ð& � ��)a��<m��VFT/�����������i��I}�`-������܍=~��@a����ϑ^��ʕiJ<�C9�� ߰�,���͏�hd7"����BY��|v��xOX�!�w=����R�it%=�dw�İwd~W,���ߐ�KYnA�[���rj�������3ǅ7���t�g�C� %�_���f����>�
���A
ƺ���1�a����������J�����Xܗe��!4h?j\���3vֿ�}��R���+�L�<X�D(J,Q[�;9���P���o]������f�����/�O�1ᆛh'�9Y�hEtI�S�*���Fsߩ
�ν�;�vOd�`����I�n���]!s\����B/r�L�l;��>��Y�k})�ܻD����w=����~�9�b|}�>Tn!8�3n��F��k`��蟺���4x�̈́/�*��7�:ê��l�9�n�l��,��>���d[L^����5��&"$5��C����+e�Z�Z�N�ж�h���T� �!�� �C�o&��V��$��yϥ���\e��v��]��#���0~���e�ڂA\��7�_ېCC5�u���1���v�̜�{E���Sx��Q�hB%y�U��!%p�n�������5X�Iwoq��H��TuJ:F��_��	pKb�^"�z#�\m<��O��$u��_=�%	0z?X�o��rp�P���IjD�#�p)�j��#�޶��J�ʞ;܏�b��_
�<LkO�a^��i��ۮ�6�����"��D0#
�%�����RA�d�1QiO�F�q�9�� �������
|�B>Y!�ƾ�b�]6U=:��7�)\o�eL�=(@Q�e͕�q=��-إ;���L������N2��z6y.��K��9�2�7�����A�q��&`�LCїW�g����Mf0ɹ�#{��Z馳}��E�=�0���ww�<����a.]�Ted��J��l��to^3ہ���K�.�"�w-�a��t'�"/) �\yм�����~o�4�B�i���{U�8���T+Ч�(H��M��Z����̹�����j`j�T��xe �P�#1�G������t�0���	�l=��Umc�	|a:��2�ʄ3��祫`��fؠ��_�~E�^������vO���GWL���=�
��Z^M���:[|���H~���֣��6�3��'1%$G�a��7���*���2㐕GV�F()����~U������-�g��P�mԓ�?"��ᓠf���cz�
��/�� <�Q���ieMa+ Ag@#�{�'���������khP[VO�1>5;i�K����O���\�6����e9��U�u~�!]��'���d���2x��ၛe��?U������)l|U����mυ��`[�,�W>'�f����A�GC���C{�4�@��O�dV���=�����,]+֮q)Λ����B�T�E�
�vqB�$A�6��Ub.����}x8�vZ�5|�/�q��+N�mP�(����'�}���8D���p)���^�b�=����������q�5x|�f�˵Ⱥjo��U��0)9�|[ ��y#������ͣ�K�-�w�XnRQ�­����-�	�U�a��3?lvequ�]�����E����h
 �t_�C��ʖ��Dz�v��,U�a��L�X�ZC���l��R�A��ǵ%�C�8�6��*D���+�o��ߤw��Qts�̓���f�/<�_b�r�͛�`:#-F�˻����
�����Y��e�_��ѝm���9 <��'��)�����[r��n��C�P�������)�V���WC���Ԣ�}k�κ7�A��ZhX��a����oEA2��Uq�/�9�9�������G��5Zc�1�S��{��=�ѽX�:��+� V��t.� �+�oV�V�VՔg��1n�
��jjh\��a�#p�=��ʵ~We���Ғ����7���'\ĉ@��KA9�Y�|%J�5^�53Il��{�${�]�A�q�Ӊ��yc��Tkpkǐ��tu['�D���]�Rbs
�d���O��ֽ��
�q����?�{n��Mɪ�QnA6�{4��t���
M�@�Q�s�zy����g���[���'�o�$�E�I��c��N�xhL����n�s��ǎ�'۠Ã@�p���s����\}-�	�M�Pc��;?ut6q��"��>׾d�ģ�kxSc��=�'���D?_�/9.��P��=�}D�������q<_��q��\H��a>A�M
��(�&���|+���"����KB$v�K�q$�K��6�w��{�l��i�?��1�K��0��>>��@Q#���𦁬�M��-|�1�6�q�RN�1;`ev���+I�$'���8G����c2e������,ntL+"ɴٶ����x�=�q�J���_�A�H�~��vYE�97���P�����ou�u��^9*�$����!���m��lpٯA��*���R�A�;e�ﹱ���<G���!�0N;r�xi��E2����;��.e	�
����Ȇ,��
�Z8d�����i^�@����fp�[j�v��D*sRB��i>�*8O�yh���Y��m)�Bj�֧*1R����������� �@y� }ʪQ�/J�d4��u���j)s^���h>, 1/��oK�
4��ξ)C�y�-7�^�����%����gk������S�)����6�.jY�`*O;9U�5��"o��% ��.�	�<�k�6o�ր>�I��}9�O.���H��f��ȡy��в��Ƴf�v қ�pؤIW���a��s�Ӷ9p��]���H�jUk�f'B'���"A��wG�<���ٔ���~�ѹ\.�9QE�1s�K��!��:��4A��j����<��f�=�N&�j��i��P̜T0�®<��$.a_��U1�؟��bR�6-LbD�B�"5�~�L[�]��c�O@�	�O�X�{3����q�|>����o�o�l4�BT9Ӟ�΅ޯ3hm���@͎)��)}f
������R@��_���� �jB-�j�:MQ	1�
��e�m�4MX`l��Ʒ{�X!����^�t�� B�2�S���Z ��g�����4�c����g�$W8Gl��,���X������ya�~s�;�Z��.�.����MDJz�U#�<.1�^��縷{{��@�����W�!��G�y"��8���~�tt���1R_����Q��l�)�N�m��3�v_�';�uM�������Ӽ��B!�d��l���^J�
+�z㳊����%��<�G6�VJQ���6�:�.G`�\)و���)�`���+�WɎ��\�%t&՟+!o3(��8�Ӭ��J=y
��w~#:��1�O'��jM�*��H���NS���I�]�ʨu��
�$tz$�GU\�}.ݥEV�7��ZT�r����}���xy�B݁�3�NXe��c��%�-�������%�v����;n�!�Ya9�������]˦����ZO��*��XR.^MX���QX��N���N��1ںV�Kh�H������ԇ�$ͫ�4<>�*J#Hi�F��E>�	]��Z���8�&����?vȢn��;M����O:}>�9�/	O�:�(ƨtjl��-\���,�^��v�}#olzH�{Y��%l��z��y�x.�%�*��3�W�{\?���X'�Hq0���{z(__���18�8GnC^s5%B� t�kV��80��9	��3:��/��y��a�E�@��A���br�F��]�.Xp�9E�?�Ɯ8wi�um���s��J�5B5ļtN�S��8���l�=�3KOn*���fl�ۆ��^�[��&=�>֣�~�gS�l�3ӏ�x���z�<�ty{�N��x��b�0�M���f�'��qy(��?���GȽ�*s�ڝ��U���52�� �+8��"1�f �Pg��]Y� ٓ�e.�O��	B,5�1�I��)n�
X��h��K!^N�x����x�Zb�H�-�Ğ\y�-tK�DdtعZ���"�0�G="p�L���.Қ��%��F� �ʈ/$&���X��2cN�~A짝�g������Q����zUO�Y�j�P4\#g�3k��]��AB$��y��uu�g�p��yo�q��Rb�a1�(���i��ֲ	��o�o�.�t��*q�\@ wb������Q�jk�,#U	�P���e��1�������g�%���WDZh &��a�9���G�R9nn��=�n2�Ŏ[.�8@p����9qu�h�x���Έ1n���=XWTX�E�cۂœ/o�~�|i������nÅ|��^v~���Dm��Oh�)��t�/���'�0جW_�9�*��|St#��2.<�	ԉ�st�����A@�dz��c�qF�)�xJ
ӕ��5�8�<�,?�>���^���ʺ�=�{��q�0�y�u�b���z9Kѳ�7D��mBP����m�P���iS���PvS�G��\y�i���
yY/X5���oߟE�A^��xG���E!�G�)Q�5� /:�|K��"z{�K�k��u�ke�g�D�Ry�Z�{�Kt�o�ybz�Z���EC���7�^�ז����n`�%d)҅2��u�	�m�#�^�<��S30�*�p|���G�@���Z���<��8n���s�|Ӑ?���!wca�O0�Zt=��߭��ހ��7��6_�~�`1���O�����Ϙ�,[���n߉Z�3y#N�w'��;T���HV��'<P��0<�������(B��a��_-�0�B����U��g��$,��/��|�u���N�,���X�$3�i��E�N�t�~��G?e�f�7�p�N�VBD#�p0hS�[���s�u��3J��(��ȫc�!uy!�7�0tS���õ��p�� #嚨������~Ϩ#=�,�:��~631�hyj{k_����>��`�I�#�l���[�)V4&�j�`.����;��v�����o�t�뱷�h����,���D��ѴLv� <�|'^tfY�n��<m:,}����m����	��pC[���ƽ���<[�z_�a��b�O0[�S��(L��f��u�����Q`B6P�Ȭ�����t���F�:ؒUY� q�h��i[�U��܀��6&����"�`�rm'�.~���m����[���2����ɇ��<���]1%ƚK�Ƽ��c����F7��I�ң�j��I���+�]�Z	�B�`[���,T*U��D��n�L^),79;�`���&�!�ǀ�Z��ږ�>����~J�����F�\{��A�b�s�b؂�e�H��>b��B���DmIE8CxѮ\��'؉}��g�l7�3�E�Y��i1��Z+%�e[�����rZy.v�O�aݡ�;�n�%0`�з#(�9�u7aI�b\� �ّ�������b��=	�e!K2�������ƈc�g�r�c��}����i@]�Ă貄��N��%��KVv�AFx�X�3xc3��Н�E8����Km���戃&�B��XckU�pXH�Ul�Tl�I�#��;Һ ��m��-���K�<K��+ÃV"��{���1�e�c(^!FY�w�2-�&�e҆��L��k�Y ]��n���;�<,P����64��gj��_�u�����P�0uvw5	���R��*��ЀvI�(v�I���dJM9(�^�]�Ff�,΅�:LSt4�B�
M�%N2h���8\e���NrF6�<�``����϶lɦZ5�9�[߭^6+��g�5n�&??~�%x)
�k��w�ݿ�0J�cKz��/��_�|	G�3�~��Bmw�V�wt��?,vYY�4YF���Z��RV����H��`AWA��BF���Ѷ��,6�hU�(����S�移���Sd���>��M�]��k7+0T_F;(�,D"���/E�%���?񀨍^��