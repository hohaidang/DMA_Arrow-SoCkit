��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛������#O��v�,�+�v���4�ۢ��䐵I����ZG;�uwUhﺜ�i'��w�	�G�1�fV�7�ϊ�Ó���8�C4��=�҇k�M��9�Q����Ǟ�H� �a�C�����c�&�|�ۣ"�6����=a�BT7�](���~�՜�l�ܞ&�f:XΕ�B�:�,=��Q9{Våi��}Q(:&o`�G�5�e^�5���3�n���� �c��1!Hz�'�<~23��`Დ�ԉ�.��=Cx�Sg����i%L�Ko΢+fC�1�[q��>�C7����S�g!� ��N�=�`�J���+].�D-�6��2�L�$\�<�d� J2��+o�nka�@�UZ�����`?k�}���m)GB�-�sԀN���9q�8@�P���*��x����4�����{�:�{�GEn?z2���zS
�NG�!�)S�J�2����k���^��I��a=��̥��z���y��0'�I�~D�l��k�5\����"ܩ:������I#2��j����P)�:{O������۸h�M��2CP+4���^��e��u�r��gpY,�o��>�CshY'.Z�C�/����;����TUQ���RF��}�I`��Ԋ�D�^��zc��,�V>�n�̤w��͏�0 �!@�1_7�VCh�g�n-�q�b��Ҝ��4s'PK��h?#�H��OqA����q���nm��<�$�Dx?1|�@�Ka�H&����w���
�tݿt��n��,�yX��Y��k������F��@�&p֤�/�QL�1~ۉ�g�y/��A�'��MUY�w�0Bb��ss>��]<��Z�b]�����<�]����S�Ѡ�EN��N:.>�U�Y~�Qm��5H�Q�ѡ`�֜��+�"��[� R���ŗnY��kek�o���$U������U+���fÊ��}/B�L��1��9�J��l��u�pU�Z��X%�|W3�_<���"`�7�A���w��a$2|�!�R,�k��か��.���E�H��㍰�P m� u$���~
�u�F�����á�ڋ%|ҳ�b}����/�t��*�������ig�����N�~֨�����=�@�D_�=��j���i�IFU�������ş������8VQ�[�`���DR>����u/�5fF���9��6������$�l>^�vV�̟�"_1����0���=�����g�o4�Ȇ��i�r&�A�{
9h�bc�dӈs��P��ډ�q5�ul�*h��`�If���f���4��<!�cCC*�<*�ʿ�"!�dW�8�N�FM@���$���歑Gۡ�47��.l���9�At�su���H>VX(| ]A��Z<��<<9i�zyw�T �<���C�]��
�� �������z�ѻ"ɝ ���hTi�D/��f�E̈�h��Kt*�ū�$:@��`���^�� ��JȘ,��o���\"���a���7���K��~~�M�1?���`n{�:a\�n��H\�����U��Yg�5,�j��`R����ۛk�@�x�G��һ��j�Y#c��7Λ�&�Q �&K+�b^�_��j������� q/6��5Ҹα/I�~�L�D�~�:��h�ڒ}Ø,���SoU�q�*�N$*�n��v;����c]���z�!��5K,F�m�2�;�_��O>����A8�� 0��+dj��<�k�~w��f�0���U��y�P�Z�6��f;N���a��?���9ޣ�M&v[L�0�R�",�2�,�i�b���`k��'�W�S�J+Owv7���)��Od�4Z7�����e���x�v�O{��c�F����V�[�lH�e�P��������	�[�o�8r�-0����9��˯�R��c/Υ�t���i+����f>�����3���)��Э�Jp&l�$:��72�$�)*��1{�>@���x��k��keBN�7.���4>wht��L� ��(��j��j��OR8{�T��f�����V|��	�C��t����;{�Ȯ�9�	�z����MT���
"}�=�����O��݃�܀^�b��=2�~�߄	��y��O���_�ut|�����$A(/��F;^U�Յ �_��Ԏ�*���&��q�<�psȅ�N$�_@hâ�
��=�N,q ��C�f��,�ǣ�?�5�:}$W�j��3��3��C�6+㍈�Nh�x��y��+϶�<�ӗ�,���o�l�;�u�C���]� �e$�Iupz��!��q�N�(m��䪚�{�	�?kc����G�ā��Vu%�Ի�X��JU���6���:{���o���s߈�:� ���Wk�z��iK��l�r]��1��� �I}7\- A�c�y�_D�[Lrv�>��?�����o��H��K�|l��n�V,)���Z�\��Ӿ�.#���{�����5�W����ǐ���2�3���E�]��u%}��:l:|�=:�*^i��?�<��H�b̈́gN�8ݏ���~4��%��0�D~p;!F��5�U(������8���av�𕙡m'1Qd@ط%�G"�Z�\�l#≨\r-�Y�x��{}jT����9Otd¤���H���N9��7'�^��\����Yh��]��>�5����P����Ϟ�s�Vq�mR�x�D�>9t�ǰ��_�{�Ly��@��#L��VZ�?��  26�VrϚ�>����`���:����#����B䄫W�'��|�k�� ��,C~�a��J���ܘY�5�qx���]�̻��k��s!ti큳#�/�S�7�]��D.����Ч�'w<�j5;�]U�Ʒ�_��`�o���>�c��X�$�K�m��vO�nǡ��I�o���]ԅ@�aq���SaA�Ǡ�L��(~�}=�y��)u��4�����`��	l�n7:k>�������ε�<������X�+���+�+/���]�
�}��y-�n� Y��$��/�"�,�P����H�-�b���>�E��|�Hx���}��t��B���Nhw�h����Ǭs0a�<�	��np���`�;$�9w}�O0�bXn���?CEZ�7��v��s��ᅛ���x�bٟ����*a�n�u���k��-�T(ٟ��we0��4�]��<�?�6��ԲJ)�o3^�j\�!P���WM;��T�*,�Yk���BG�w��l<:uZ�|a�J+3M'{�7�٣.����jo�J�DN]|
|��V+ȝ(�hP �?�.V�'#vس>kz�h�5w�|nk�����s����j�U��
�3�%b�ט��Fu���(o����xH|F�C�I-=��WY}1MxW���r,�V�M�Mĕ� ��	ҩ�@�����ض^#�X��kRۀox�n	~_����L9��u����n���fޛ�!�l�uS����rc��PW��D]b��<O0XQX�*�LZ3(����m�����]J?N�����`+�G�Q��0��|����@vo���� ��������t�i���
.�:�x�I���Ak�ַE�k$-�-g/J<�Ѱ�.�,�H�W��+��8���w	�����'�q�xV���
�4H��c�.�}�`B����.f� <��lp�)YS��L��G
A	��w�/h����\�m���P|��[;⡞��
2��'U� O%	<�c-�f!�g�/�o��	�0��MI痥� -s��G�B2�9�Z��sb�q���&�tt�<��8[8����Kw��1���n�SW<���Mъ}�����v&5�G��������8fF�t���i�-+�o��]l�8&rE:?�r�K)�s�|�%2�Ùs���Oz˻�[�rZn��0~[� �����CỘ�6���Z��9�6�D蠯qo8aMx�2`�����z+δA�|`Qb��l�bj�:��iMEC(@��x��UHl�_l���u�TgV�nOw��~aryXGt�k[ pEGtf��Xb:{)#/���� q�r{c����^�����\��Q��S��R�>Ii*&��8M[�߰ 2M]�ln����t�����҇��;�0Y�GY�%�϶H��6^����˙ �j76^#u�f��:���1��|��ki���}j���o������;������O�I"��uE��_'��zQ�;S�S�Nwۇ�q��͔�g�03YH���5���������DK�V���馱�J`��u^| �T��_F!���O�lG[�":�gT���S�Y?�
��89�̔[��].p��W.��,yAZ�\b���UJn��e�S �Z)Ϳ��7�:�~���Y�	�^��2+�y���K2�`�f51�eaټ�@���uR�ʞ輢�eZ�(;A��->�"0h/�6��t����J���X�B���.�_hi�F�����Ɏ�L]��ȍ�Vq
�(����]���@���fw&+	����*U�X���Q۬ O6�*֫�S{Ҥ�M�ǖ[Z��Q����FR��'H2R��?�&l�Q!��<�!O�}��S�w-�T�'xh��F,��Q��i��i�o��V��z�Pր�E�4��?���|�]Q��i_�ԭ<Z����c"��Taz$(t^ ��#������-�+����I�����V� �*�U�p��wm,��t�(��-�j���1Ko���;%ԓ��WJ�(��De�O�o-��J�u�Iv��]653[��aqm�m��*�QN9�~�R�f ��(� Z��%�ˆ���#��w�7-�ے����WTCh�i-T�.�P
0�=�"H޴Q�`Ph�?H>y���,�w���z��L��E�;��(�i]j���UM�n'3U�G�G�p�9Ƿ�:�ozAƇf=P����dZբL�Fhh@�>f��n9[�CM����i5J�I�ޒ�W	s�؇ѱdD�R.X.\���^g��k(��[�[�oZ�j����RCr���������S��Bhv{{n��V+�&�
tȅS�X�n�II=���ɑךb�N�C�K�W^ϓЭ\,�[�lʅ�KQ����bʆ�&,g།+�H#�p��L��o��X�z,&�v�c^_�M���}|��� {�å�bMߞ��K�Cƥ��G�
���L{����_�<�p�����g�zn=��d�/�T��wlc�ڕ��p�P-|�l�5w�����q�v���9)O�U;xh=��D�鶽����ʣ:���}"���({=�G�HH��+d�4�e� ��o���>B�o���:�'�-^��-+n3c~�*�w:��<@2������s5�~�0��_K��p�8r=�Qk��7���v�����������2���s�5L:'Y���(
8�3N��h<Q��s��v�]�N�`�y\��*��rm��j�iu�>3|",�������������A*Y?�2�*�2AY}�Ԍ#�A�b��j.�z'R�yd6IJg��ĉtCS��X�b� �A@���
��!'�6�K�Ї-�1Y��?�����/kpe�ϴ����ۃ�%DS�I�h�k �ZʚW
`�Ĭ�b�O�ё���MRњ.���^�f�3̚_*���K�� Ϊ�	�v�=ڈ��0_7�O�D������.���
�� #�D"��S�7`���a��u�3�.�d�J��qj��t�TZ��#=I�eZ�L�%��4�U�:�b\J Ėy"��'
�ˤ��PC�O�M�I(�Y�4��'�K0E&�KzB���jU�CeL�*3��E:i�����@4#5� �X,j�Q�6��Qe�oۺ�ԊS�PQE_��\����9q+FW�2��F����R�h�n��W\:�q�]����=�h�L��N���P���D,��([����R�OL�5uM`E6-��\�$��h���Hf��C�OAi�NЙW8�!Y����F�(���Ap1Yj*
��r6�JJ�i�UX��S�w^:εٖAzGTk0�!��3���(�ئ��@��h��{0�f��H!�A>��v/-ִA���̋�8$}�zX,Rp7 ���h�m8Li���s����<M�`T�Z��ȏı�(s����&��Y(.ؕ��4��	{�3�10�����@2xQ�����:K��P�G���n�P�A��k2�Dlq��l���Q� �Ŏ�CFr��:���<��r�:�}�J̰ɼaX�����3�
��Ɯ�j��~�
<����=��W�B^���p��(B�au{>�����bF�a�t�/'���O~^�͍�1w���I8�3@���en�3N���m_����E���ҧ��	���"|��P.�O�􆟿Y(��)�0ձ�w�����y�iW���ݪ;�:Kզ�1;�޳��:���˒ ���`?��h�x����y�~\E^A8��T,�.���`(��P��ѿ�,����Q7j������A�{�/����n@t��3�`��D�D����5[%�}�.��`Ǖ���U�E�˼�۴��fN	�:�1L˜�|Ln^M_��������󅄼��f}�P��B
)�-$����F�7����%^.�1n��T�[�*�-Oʸ��(�C����'.�U���!	��_cEG|˂3��0A#M���gD陪r!&��3��Û}���l�����ۊǽ�{SFx3֣Cr��b��W��Q���0��@X��$z���7�4m�K�mM��%�Y�G)���sL|>�	�v��n��DO0}�b��E-�I1����^�����9��kptĕ�"�l� ]ت��|��RG���HK������+����dGk��Q���O���s�n0����)��z���0UvfYv0Y�^ܗ��PW�Y�?�������Z<�%"�+���︶8�F&9<v�B�k���٣^���h}�����+A=Y��}r���u��8н�4��rp�R�s!2�̲�h�@&1d;�1��SUR����<ib�{PCu��WT�4�Fiq�09Q �ٴ0ھ���w<���N$�쯘8%�rC3{Xo:|:�N��
�!*�τNP ֮���V#���n(�}�� S�R(;6n'M�Q|��1zS̔/2�{��ڨ��j�d�4��+ÓR�Ɨⴟ�%s��d�0�ohR���i+��}4w��C�xR�ͭ�#�'A6�K!�����bw��v�~;Z���I�8W����\� �nM��.�T�/���-~��p�� �T�<���"�'���K��5E���֊^�����������w��&Xor���I�l*6˻���9D.�,��[����E�5�m�Oގɍ�C���P���b�А�5r$V�Rl���_�����g��,,Z�L�w�O��Я�pEQ$�x�+de���"�z����H�&���c��6������u��p|н�p��Gt�c(T��C�XI�E���a&O}sow�TP �PQ�c�Ņl�=��ނ�|-�25{�gM���Y�������,N�B�'�4݂"D���g6nv�9X�zC /k��h�	�g�o�Jp �{�́V]�W2�,X���"��� ���?���_;F���,��tBU�&6��Gn�9S81��'��h�>Mʅs[�bY�H����ac	�.����md(����"mp9a��M�S�3�pg%̢�e�/7�1~H�tL�W�:��G_u߻*����"B(�N�8�y����T{S�1|��l�z3�V䊻�#׹x�V֕�����/`p��.����ٸ|3��`z���]b�z4���m�TG^��z�/vx�@0�޲�q��$,�_R)J���6egm���b�Y�QL��;��rp��FV����F��QhD����qn>�,�>hlC�SD¥-�=Y�ɏ��)�,�U(�p�U�3�󍽲kS��Ǎ� auru�g8�霘q��(� 
�F/�M����=,������ux	į�=%�_TWQ���r���W�{'�L|��uw �`n>���!l������eMw�b��s�,��|Ψr��Q��P!�er4ft�H�B��Ź�~�L��y?�P}v��'�@�M����y�bgx�0�*aI��q�\d%���5Y�����"{2
��=�X�5z�;���Ph�s�g���2 �"y���`�	4o3�E�V��zx���F(Z?nm�z��vGv�'$0�� Ù��<��ܗ	���9����OSBg�!�̶s@I�yOC�yY��G�m#�[� �Nk�tK�l��Z(�[���%!�*q������	� s_-�� (JM��8,.��ݷw��m'3����E���2��b�Vj�����-nM<�k���IH'��ެ«d`��(0�=�jf�|!��غ�� ��zN!7m���gb�|�]���pۖi��6�Lp�/�@xgb����c�k���-��i����/q����X&�ʹ�y���f}�B�-d/��G��Y�͔h�_}?��Z���u:�U�+��e֟��.�*é���̱���VV�t�>3 fs�9��]� j�	 J� �H��%��y�?z��d�ܣN'�z��V�9�~��J�E�DXr-�/8c������h���%8�B`�c��6�l6W$&7ȘdP�`x���R�	����s؂Z�FU��~ UM��"�ty�˭��r��}<]GE឵D�f%R:��		m�����24���F��6��4Q���dW޷��`9�Y��qi�ߋN�h�$ɗ��M�'�'��DY������ORkz�(/���}\JO���l��E�MY���(�� A���R��:�/��X�3H��@7�����
n�ڟ�	&S����S�ɨ�ς��+�l&}s#��܀c%������7��_g�Xs��Z���r�E�ճ*<jV��c0TҪQ��_X�ߥ�0(�v_/Vk��7�ց���`�`�Q}}X'T�O����~�eg��C��hf)��4��">v`yQ�Jç,�󸑾� +�����xv��
���XQ<��g��nt��]:����w�j1�`��8O��D@���3�ƯHt1��p���v�ܒ�Q (7qc��m1E�6�3�c+��
�"ґ������Srtu��&����󨘚q��\���y˅$�K�tv-�V�J�
����^зP���#ؑ��sW?zYm0�{(_������:�^���8P=.f��au�p4������H"�:B�ʓ�ͪ]�dB� �K~�b�դ�j\�N���$�< |�m�*d-���sil	�c��k.L�1��7�dk���㠳��>t֍��ЧO=g�3 M�^�,{���Q��&٬��t,9�h�[���4'�����C�?���4�P׿��j��"�H���ʐ-�/���P��
5w~t�ou��Vy��`%��W6���#\���k�=+���X2���nt�oTd,��l�0ˍ��鋛Ի2�i�&zh���鿅�W<�v�0S�6�.&zó"JaΒF���%߭E �&4��^����]�v���wŇ��d�.���|'T��.����,?�]�!��x�4�.�/.A!�� 6�0���Q"�-���>���_E��A3A�r>��|�����**���A2w"����`�q����噤���6��	{�����	�m���c�G'5:S\Ҩ�7�˸Hx��p�K��Ӑ�KiXn���zRZ���:�{��v�^���%w߱��A}q���=?yD��g��ւ�C��䜐xјey����ىE�&�m���+X�Y&���>� c�}ǇJx�����[QnA�����w��i���ר��T��s�]f����#�X�h��
�I:6��L��#��V`�KχƩ�I�RP�����J�����Z� ��O\����Zx��0Up18�R������z=&R�����7�6=Ĥ��|@X��Rr���u4��U��>���(���`�x����K���OĂ�Y��l���ɟ�>��T9�?0�gΓ�AJ/P2rZ�\�Ά�薊��ݮ�p[��U�O��_�Z��);a���!D��Z�
8�!��G�~����!�+�>O�jO(�x�D]�])R�	q�h��[G��R�-)N#�)��=MR������c�^��m0���Gx0�).�XKb�H�?D�Wr۝�j��Þa%������Kw�`��[��#��h�����d��M��k^Axx1�:>�
�.�e�`5���=�
�b_^�6s�j|���y���K�������j鴔d)��0 g:����|2�ɕ�R:�;1I������� �V�?���9�&�C�Gld��Z�����
g�̆�+��JI�"�,�s�ո/����@zB�� l�9�E$nq񱷋�U����6�aޛ=�@��7�F	�Z!��{�4T� �F�9�;�u5+�|s%^�HJ����la4��.X�6*c�W�  y�*�Z_�֣Yt���Ha,��'�_y4�G1��B��oN����XuA�>�y6E�Ic����4�b3� ���nˈq�J�����+��u��'�5�\1}��I��P�m7O�9M�O�p����9z���;a2�7�&
���b��j��O�e/��ũ������j�F>��� o�B����b%����[*�C��!��$��Q䴏J�+��>w�5�Ow��;	�'����r���= ��]� i	-ʯ��2��ũe���(�N�
u)�T�Z��Y)^o���ѥ]ll����u���"Ą���_��4�cP���%Yˇ
�������^a�f�n-b�A�1+m��ٟ�jx�͎:Á@gWdty�\�e�d�e�L�V{���s9��H�n �g&�/	��qy2ݏ��z�,�n�W��ړ�VC�F2�yp^c�+�"�t?X�"n&m\Ȇ1��z5�V[iIB�x�<� ��R�.Ƴ�(�fMS&�F���IJ{�dGR�lw�611��6��<��Ո�k:����r�9�\���>�ҵ&ĮR[�-U����M��k+w#��+��j��U*$&g\tJ��]��̝��#����e/Z48���&rA��Q��ū2��KX��l��\G"���TMl��N�8N��b��ж�&��;���Go���%bE}`MK�^���;X5e8	ڈ��T�Nm���lx��B)�}��̓�J-�?1ߑ�5���}�;���?�*�l���JO�� �&��i��u��2G�Xru;{g����s'�,Xui�=�_�68d�7Q�o���P�1*��Kv�X��ϧ�C��c��֞���j��șk��{��+�Nzl��������i���>��10x�1s�|�b6���!~r����T٘�~�0�������6�\&��7�lH�S��K����.���0_����
�|���9i�nHٮ��(�~:�+�j����S����Y��r#�a�Q��@#|������w
�~�$/���|�@Y3���������X���J>	�\v`�o9�@d�Pp�M2�l�ѷ�.?�{���#B��G0 ��a�fC}׽��<)��t���5�57��T���E���+.k��#78f��ڋb�9@�a%T�s i�qa��Vb��Ӥ��q*��DU�⩴��}nގ@I�&��ֱF_ݽ���\�*�Eu?�]�x;̘k�,t�n�^����T�~��W�p|���sɪGh�K
ǩ=��l|:`U�V
�W����~Oκ��RWԹ|�����R�_> �����ϒ�0���X��n�\��q���Yr��'(?=~ƾ"t�쑂s�,H���bBB���g�vy�@?c����'�А��fIm m. r,�n�`$�%�s�e�9I1�n��=��G�4�&	���7�
���eU�~�ü���b�(��K������G�Q��*Hf-/U����m�W�I%NtE�w��8MY���ޅH���x�ju ��,���Ao�"C_%���1C�^}X0T�9��ZM6�P�lw#O��!&4�htmh ���I���QT]E�p'��[Ό���ΙD��0a��7����A�|�3�������!��.ioѓp��ʭ�×��hn���X��&��>�#���z)fKR������*e�k7�u�Ҹ�X���YN>(��=n�q�\�vd/Z��H�P������.�a����Y����:,#�����ǰ�j���-��tjh,�PȒN�?R�	�R��; �4����;j��)��YR|���B��ĳ��x��ᇟ���k1�s��M�*m]Xo�Z���UP���&9��2�@�[W<�[L5�x"�c
�߽Xn':,���y�ii�hM&��_|$7�FsGV�l��C�}\�	�
��[�PCY�q��[�|q��D}Шp�[�u�U�2��ҝ��Z��I������ (�����U�����T�з��a��7*_bGGI�wP�n��3��ş�ŵ���a�����������Y.�����A���ZMD�ig�}�/k��4�}�A�_�f�I�XT���߫a���L�\�=�-�E��8a�t_���Ix�L^-q qc���j��Jo����yՠyۈ\�Or�+!��%��J����q0�Z��2����(�xTR��1Nي+"]�m�lT!0�3�n?�#��
��ܜ����{�P�()�u��3p�"�{�U��Gm)g����`3�%��Ď�C�ְvC�o��U���aQ�(���m+PB�!���Dv<�>�F��K����k�R��")΢9�^?
Er6�!B,ɂ>�)r\3&�؍��ZV���*��`�7��.-�3O(cM���df}�A�VA���,���v�u8���`�5Y&5���cv����g�,p�h��g�vU{��(h�r�@��_��ʪHv�eVç����%Lw��NO�@�I#�O��f�)�93]����p!Gc���Jr؝n�Ԕ� ��Y��{�Dv�"=�}J$O�]*��p'O�[�xF6h
���UY�Pu�c��B�S`n]��x`aD������p.d���ݽ���:HĠ�x�i�R�[�\�Ȳ��~<����Gy3fG!��[����ӢIa�D!���|a�!�Z�s��k���B�C�d�
�ٙ�ZB9�|�H zX�O 9+TU�k�����S�Ȫ%�e��b����I�1ܖZL�F����$i�4�h�yJ(�]+�e7{���Cl!��	gU�2�Fь�P=7����F߯����g�?2D��=��$`+=g�\��
���G_����k���h�:5��<����n8���;�Y=fY�xf����6�x{�EF���c{�����{�B�~2��ם�� ];����� w�va�*��z��ڗ��f�f�����~̊.�3���՜�cfw�@	�"f-��,�,J������I�s�j2���,&���S���Aa�6�~Me>8�CY�7P�۳��.33��î@�T�2_�?`�;Iǽ;�u���ROz_X�������z�Vi..�]�3����������|{�$Z�z0��MW�[ '�U�4ض&�jq���C7���H�����y��#Ygi��G�d N�� ���1ea�1?�_���^�E2��oL܀|�PN<����������cG<��-�O�Þ���A&�[�����U�8���V\��qF־�]Q�J5�
�č�}��&��K+#��_��� �u��Sb 5�]��O���mIU>%B��*%��I#^	�S����Do�u��ܝ��5�a����JC�-�rA�y�J:����}�vѺg���H��y�S0��2^�`���'���~Zŭ+չ9D�b�18d�`B�7Wb��̪����;�"4�}mR0�p5��aΗۀ����k!q�=Y p1&5�������Eg��WB��Y엙م� ��aF%T)��h�
 jU��i�`Y�	#f��i�vB��9�  ��#��b\f4.$/@��3�ͳ�O��Ȯ�X�+T�����&>�#Z��OX�Z�i�����@�y�g��S�>�=�=8��l��N�H/A�����6?ՁV�̘�,e_���x���b�8��_t�GS�Y3�T+����p\��!�#}�K9#�J!b&��:k9���@@�j��c�ٌN�K������D^�=ܳ[����_4S���%�-��
�,jؔ�
�(V��-��0����n�5�l��W�bá3�����Ҡ�{� a[*��m��6v 3�c�by/\��?8P��(���������
����ykO�ٽ"YC 8���x s@m�K�,W���4���,eZ��Ʃq�ȿ�YM���s'zN��3'�?����uc�(`��J���u1gu~�򨡸��t�8���[++.7LR����_~6�6:v��'�*��BqddG�|c�VO�W��*�H��`��۽�<D$��}-t����v"ٹ��8�ɝ�� �d����m>D�_�����p��]�x����oYs^G8�Mm�wI����x}��/6B�_	�Gk$����E��w���Ɗ�s����sp�
X����*�E���b/yu7:�3��>�Z��NILDω���w���A�V����������ß���P4���B�awS�o���E���)�G�'�pdM��\+Z�ƕT{W?Ż�vPa��n3|LU�����ɌǼ���p�Ui�G������tQe��8�3���e�o�c��f��O��Y��i���P�ʄ����ۡ�ur^�S���Ӓ���-�Ƕ0�Ur\'x=��4crL���3O9��&H���֪��`,'�g[/X�9�}��A�8S�����Cgh�8����/ڭ;��5��>?�)r��h�����t;�f�8,hh��ֹŋg�?�\6����QMF���uB�������;�n��cU��-�A�τ�;F�{��?zB�2�_�0�if��It@��*�|֊�x��^��3��8��5&�� G9u	B7���
�K�f̃rN_t���'0<��a�X%;Ki�B2�`��=�G��]q^A��V�0�n���k'� RU�mH<v�U�O~~᳈��8�l���*O�r4�LL���� ��q$τ�[��EYj�	̉�{�N�U�[aިB���q^E�m��(���׽�?%��d8����}��].���z�Ǘ��_�Ϥz9AU�Y�b��o���������J!�fb�#ڿWz��<+�����֜���}�.�Q�@�E�:�g��F�.d͓�U�#xwx(�_���Q�����m�Y6���s��:��x~ZɁi�?��$���D�ő�S����������"T'�p_�&�������w7o�oПY�[�����TĿ�K__p@D�ܨ#UneX3�ǵ~��R|-B�&�s�g.�gұ��=�wz�@K/�W������q�>��ƌ���æ�����,�5���"�Jd<:������������0�$����%0�d��d��@�%<��R�m ��$�UP���I���w��Ee[�煱�z�CܗSs�OSݖl�!X��i����^�C�"��,G`��Q���� <:��%�V�c��]�����:ʽPm2S�W�߼g��(y󨸃?�(5����y&^�D����O
%h
����Z-����<)�<c�چ�e��+�ywn&@��{��fIHJ�)��W#t"F�{hL�5'��`�
a��D��������F��u�P2nA1r
�o�B���m�'�k0rꐧ���%I����b	z�Mte��&8�+���G��?�S��#͓g3Ɓ��@�X����}V�Y��]����??Խ`l�XI�0�L�E���*��(*�1+�.�\)� �5��d�r�l��R�kuqW'��S;�c]�p�繮J;)���������x�����j-�%igz���D�#g�a���h(-e�$d]�����4K�L��N�p~�# N��-�|���d�0�9A	��g��gEwT���R��5Y�gN��xqhP�|,c��=q�m�E���(iZ���:�r�i�>���O�v�F[�[�O@���o����a�L	Y�4��i���٘��:�����=�B�Ct��sI����h����K���`������!TJKX��~'#�{� �J�_��dcH�B%H�G$�J)2 &�k��#'��ᜑϦHJ�� i�老[�
P~7z�bn�s(��^R~�|�=/��^�j2����["rz��&�^b�-�}�
م%Ǻ̱M�}C�����#a]6�M�`��si�}Z=(=�c�S��q�L�����F�Z PP���.���q�w�QJA��A:-D0E�r+����z���v��	�?�J*6�� م�����f�ꠊU��/|M�٩;�3� 	��/���h<�:U���\��h�"�P��/�^h����91L����V����F�C�D���K��lS�a�XA���#k�O�l�Ć2��<(����ݮk�ځ#���R2���L8˘o��F�lb�CI��ϐ���*TZ@�(���X'?�t�;�� |���|�O��h�� ������u�:*,��K2���L���������� ��(�Z��5�B����!SMJi!6"ċ�}��J�+�m���[��b2����$��|3�i/.�S�lߝԏ@�R�1�0O��\�]Bh`�;�ag��M+
��ꕘ���v�B�sb�6�=��hJ.�����#�v��4܍�S(D�f**f�<T�t?N�l�#$��ی������b�Q�AU�;���zю���]���pJ+�yL�'de<آ���6َV�"K���?|{綏�v�CR�c֝�Gs�_:ݡt�i�}"�C�d7�%濣�Kk0a��;6S�iH���M�`����A��Y �jz��v���%Zj�.ɮ������Jj�(����ݚT\1���������⢠��R#v�f6<��5�I���^�M`�!~U�G��H��j�� �;����t��^68ADM�M�!�;����wh�Z��<WZ�3y�ozޚ;�+q ��JX �;�q|�U1˗��Y��YM�4�Azm�
c 6�S(�-�|z��{Ut�u�'8����_H����Yx��S��A$��c�ؔ������OD��T2��su�;Ӳ����ܔ�t���=�	!���$�}��͸�K�P	���z|Uhi��eX���q�K�L�@���x�>����j��U��"�r���$���N#͠Sg#��XJ�ڣ��B���FF0�r���)qΝ���z�9���BMf��qE@䴠�^{�Q��%Ds�4h��O��aq�7x�e��Kci%6ʁ�T�	���h��n|壨B�>S��`�]�
��,S�@�ڈ�I� O
��������[�P�deΎ��4�}rh�Z[�2I^f~��,�^:��\ʑ�C0W��ʰ\4��y�)��OáEnP���x[9T���s����Y�.���C"|%��	u�h�Ug�j_,�Ьm�i�g �Ȩ`������ �<�03c�?@���L�{�:�种(�8[u�4�s3[{[#;q��2�A{=>y�k�Fm�P�?%A��U�_�T����$"M۰��/{R$^�������f�v��ǭ�U4�u�1�zI���D�d|	t�n��?_/�[�Db$%Å���=	����EK�~��2"9ƭT@�&��?(�;Ş���v]ƛG�*���(b�M�e�� y�g�{��%]�&d�_���+���=�MK�l�ʚ��E�&�1�Rh\�8n>�2@8xv�B�]�-��Y|����W�~:�~���{[���lS�J��c�'eR�*b!~��遆�BY�N�4	�j��aK?d\ �U�̅��{C���}�s @�2��oՊ7�Q�A��b�,#Y�L�BD��p�k"���k3Iű�"��0bR��7J_HM�s�ž��ѣ�6:���1P�S���Ux}X�P�b����G�?��@�Zt'�m���T|b+�,�"����8�ìUv���k[�|��i��9�аW��?0]?TȠ�����F�8Z�	$�kz,Y��S��ago� I�N�;�&i�'�1�Β�� ��,(�,؜hL�烦d����[��{�>���4u�����蚈h��q*:�f��N��	S��z�C��R,�P0N���{�o�k;�M��jO��� ܖ����7�L'cJ�Y�n):�{\���_�8lX���T����,	)X�5��e��qa�{XL���h�5پ��;���ۉT�pu$5Dǝ��aJg�|�lqn_c����@d$<��uF�pou�ޗy��}C���U�8�7��g��d���?����>����w�Qܪ) ��x��O�_������p��F��,m^�&k�I'^â��*t]/�V�5Y����L�Ja�Gn⋠�����rSZ�*s�c��-M���<����!!@�5�ʋ�����ו�sr��(~��p����Q!p��y�j�z���~a���1�$oL�1�dtU��p��� ��,��
�H��1���:�R=h�k��^ǹ��cO�C�v���
pڔ�hJ��h=M�LA���&(��S��-3NՌ��ϭڼ��i�|��iٞa`�[	iۈ�����W�$�I��5�_t񚱩$c����)��i�wc]�*\D'�eY�
�Gw�1ll��-���P���H��V���"�`��d� ���Ԫ�.�Ya�2�>��|x��6%�`��^�&��%�v�+,,Û,��i#�H1���,օKw�ml��xOk���.�凅C��QRYQJ���Z򚴓8��VY���/�f�b´2�;\[��%���.�Ez@����s��l�^C��kgu�e�&W1����?��F��!�\7��f�����.�Y�Q8�$�`���I~3<"(�z�s<�4�%A_%S����}�B�_Vd�e�Ad�0;Y�\��͟�H^�@���3���<�te�N��GN���~3�іS�e�����7e�us�\C�+�k�b�Y��a��A�f{ԃ~�cd��糎L;����k��_��)�_v����L���K��L=Q���R�Wޏ�L�3�]M?�ejz�x�A@ ��b�Ճw�喦����dr���Tl;B�=ܷ��W��R�`����M��g'JN���7?*q,���vˁ>m+ �g�J�𷁐��/�a�H:�ZM/�ӣ�|��Lb��/C�L/�$�,�a�1[��E�{)1���#S�Ov�%U�>tV��i��T� ���Z���o�I�h$���ڃyJ�p�mk~��k��8��p/�y�M�b��8R6.=wA�ST�]ɹ�.���i���2p�k��{��2�O"���.��#�d�o����-eە7ڦkX��:��~�ȼ��,�h87�[��ϵ�\ۺ|M�H ����;���	�4H`�}���`�;^7[\.F��l8��d�,��]>yP�>��!���
5 7�	^�(�gh����^�a��F�O��us�s���<�U�e�j3��R s�m���:�N��+,@�����ޘ�T(�(��Z����N��;��4(=0sG#Uӻ/�|�*��|���3@��T�l�z�T���c�W|���S����V�d��nX�Tn$�[�V�[�����I��1ף���$�7I4,#s���,�{ ����/����eq�co��$�x�>���f��׵T��:��p�fQ�V���w��{K�(�l�l���P�;"0�;��2�H��ة&2�N5� MM�`O��@I6�0�oyb�V4tb�!�T����לߎ��엫ʗ�;�zr�n]������J��C��7���$�I���p�'�$����,+s�{���(��R&}]�h��u�]NF�����h��)�̵ŪV��2�{�Mqd"��H�iK�7����hG�ZB�Ɔ�϶-c��	>kj��A����J�A�t=�8J6�U���y��t`$><�\\5�k��J�*�hy3�8y1�d�\�V��D&c����`WQ��ERuA�%a�.�5�p���xO��_�6b��l�O��R��x���HV9D��dP�K��߻��$��g�ٖmn�G�o�E��	��u��ȅ��2�W�E�x� >~���Z$8�p��s#�_[b�|��5�4w|#�"��H��?:��xreD"�uG�2�qΌ&���9�=�z�{�����2���0�Hv����Iip+
�hڬ��[�P�iJ�/���
�	
=(+��q���%��ȞͲ\�8�J����䮤mB0{x.?d	E�E�^*
�}�ł�)���MY�<0Hm2h�!���1 �=�o�8����E�9��\�"9A�zX�*4���Eʘ^V �܎�M�(�+X�iO=��@J�I���v����h(��<ʟ�Ƒn�/o��z��%�!��z���r��5MB��`�'d��oC�K;y�h-��%�K&�t@T��61�ң<Ӌ�}��+�6��Z������� w������c�+ Xm��#�Sv���i����l��-��xE���5]�W��[��#�l�#��_R��q߁c��{�I\����8�w��ܪ���������?_x��oߒt=)�ׯ�5�̚W"Q�c�^ÿ�D�Ӄ��T�ݨ�2���y�j��s�W�HP��p�b�GV�q���ƥ���D�O��~7.�D�<8N5,{��f	ay�X�#��Ԥ:���ڶ�S�#���-�b�B��'��>��t�˃��V��aˠ2\���樛���$����0���
��=��������������6Y0&�D��m�@�����Y	�nQԠs�+��E����OJ^ɂ�c��-�k����Kݯ��~,12�����ϖ����u��M��TI�F�q�}],p�4�,�gz�BK� ��Ny���5�m1�1�QRy������������_����Q���rE1�䗰�M��w�T���JΊ����E6a��c �I��e�( ��=��G̓�$�a�d�U���~b�u����EGi���/���8�u���dY/`q�_���R�=�'#o��x��eG*���P�t-cuwĔ����9���&����c|�U�V:��)�ܷ;�"0�C��c ���3����:a�~Fo�_�,rm�e�� 5����IBO�?�
k�)㈬։1/a����U�)�p|> ȥ�ib,�K<@ţ�]�X0�	��c5�����IT�����6�~��ڲT���(a���������ϕJ��~��[:R�c/�k���������ˑOF9G�I;sā�FF�/-�hN��-Sl�_�!Y����)�����:$t z��G�
�xT��X�F�%}��
m�v4�4�>�n�8�r/��-=�=e�RM���#�)R�;�_��a��˟��f���=X
�s��}� ��=��`*U$�,c�"��R<_���~��/�voƐ�#U�'.M���BN���*�t�L��ý����]���|@*M�+]�efi��,���u	(
������I歈4>��daWU�4�ΏX��/D�r>g�\�K3L�؍��H�9#m@�-#���e$3.����7�u����O�K9D뒺�!���Z���X)>�d"���At�8��p �\�8�0k�D�&򤲨��Ϣ�[1�s��_(<��K?�H�QP|���R��&��o/J&�+�T�PF|�^��Ö`H�[쮴f��J�@,�D37sZ��<����b��;�^s�����J̀�L'W��V�Rl<b��x! �����$����&gգcP^rR=OZз:��[+��#ҴQQ��)A��H�j�iO:n=�u�� ����q y��ֶb��nʎ��K������M�q�F��Aڗb�S]|&�	�舣uH���M|�P�0�����l�	���0��&�s��"|� �����?C��S��+��v�M%���[�g��O�fPQt�EJ��(���:ԟ)/˭ռ����[]�F1\+��"6�Dl��Ɉ�d�9���������	�Q����pu��Q����_Q��-�r��)�D�+_���q�,i��k�-�hS0����S��B� ^�R����_���KsA�v������o�F��q&Z��`�2&��	���#����������)V⧑¦V �	*�FV�!G���\��[�KG5J��YDR�_��1����LMLc���Wjdi��Xfr�G�QH-+|�=_��<�d�uD��|�՝�w-�ꏍ��An&�ύ��r Â�z�ԓgH�`[��j���"�K|=(w5������p8�j�f�F�.%�zp�H�>}���+��(���UI��3�D�~_�~_���;��	�D{�k��U��n�[��V7��'ϋ��Ð�D��}���,��a������1����>�1�F\�!J'Ql�yHǣ�lK�	�G&��,�h7��Jz���\l+�-K��qTR@���Q�o xC��d��v�#M����a��u}	����-iI��ϕ�2sf4���*K���S!��?ꭜSz$���3�tBV�m�zT���c�q_�%�w�2LQb=x�`�#�<�E]��o7!�Q���������X���e�_�|�+-�7�vi���˕"��
�����}����������y_���leq�Ag8(���+)����p����v�.A�]Q��)����#�Ԗ�f����3��/��Ѝ{�g�H$���@\��l��t�&!��,�!����eZ�WZe��1�}���.`A:tM���F��/\�ؔ(�U>;E �M����BP�#�1&����˲��{x��bV��e:����1k�U�G"J���ZK�`W��~�6�,��CU�^�@�Ỵ) �z��2����AV��NL�'�s=�u��Z��r�+9`R�B|<߲<Z�L 3�V��3�M92p}�5��5*z����uͿ���?��(r� �X�[�VxѪP��3s���Ŵ�����I҉%]7-Z�6�;)��S�m�*��s��\��<��-k��pw��tdm�y��
d����*R�du��#��ҼL:׳��,2K�#K�I>�lʸ��[Fn���^s��Ӹک�p�шϷ��-��*X(�Q�ސ��#~F��C#̏L���Ч9��]F*��'�ُ �`l�A�C-��)�R�Y�!��&A%�UL]�!E֢RA��}�R&�rn� ��hF�HQ�TՃ!k���E��бa����O���;�$���Ї�g��e{�~,[�@�)̮�E�~Hm
<�°���+��9	}Y$�*��k��§��JQ�=��w�k�v� ������g'&k�n�W�F �����u�_�yJ��y\�H��'�8栙t'3�ٌ}��K���`P��-�K.�UJ,<�6=��Chy5f�ښ�[����Ms������裾1ߤݖ8*�||�
_�Xj���2R��۲$���ݿ�ȍ�M��WkN�NZ's%�_q��(>��
X	PW-B/���,�AS�.���
RЉ� z�^�Zo������_�*;}��1	���4�r3��(	�y%o��������gNմ��jwe���t�n�҂3J4�h$��R!�:�b��1��	յ�0��ɥ_ݬJ�w������c��쎤)[�+�+��q¶����1���Dm EDEuVm֜�;���.IHF9u�#�>���%x���ze�`����O��Z���Q�X*� Z��l��	�N1/�G������c��(�H
er,���k�&v,KS�'f������Z������$U�S3��Iw�,���!�!j5x��Cæ]mx���o+Wj���C#O%�s�i�8�t�s���������t�E�3�:M�.+;��=�3�;��1�>C���������%w�Bz���*=�zY�k��X�9b���,��ɋ8�4�?^n���0�L��������J2��2��p�e����>=��h�?�����.اJ�kMk&�d����0O	�W.�W�,���KA�h	��Anͺ�"�f�wR���9����(;]+H��Y��q�Xߛ�02��=P��z�q;o��NnG�$Т��hI�Z�*q��RA��e��9����Yz6�]�v��ZΡ��}^��8wc������ݜi���;��t��p�6tJ���Ck���������#�$��!(�C�=�W:�7ɫ�M��� ��#lZ۔���i"i�*j�y���w�<�5�C�E��(�O=އ�ST_}/W��-5AsPF�=wm��MM�f���1۩t�[�~\�@��t; ��jx�ky,`m6P*��:*TV��8fD�����/��{�NӃ�c��YysWd0X�"�\�^i�(!�-����U6"b+��-o?�<��	�U�b����%꫙����w�N��#�7N1�E)����\R�o�K��/�lT��z�M����⼜	/濈��BG�:�i����΄���`����L-2���d���{�>�>c#�X&$�m��<w�R����ܹe�
�(�5��{f�g[�t/-���(�8x\/���4ڢ��Geh�e�|d6c5h���i� R7�+�����u�F9��^�;`��7_��01s���y=��ة&M���3\܃�zU�o��7'q�����|���ڈ�k�b�jN W�4})Y���s
���ziX�D"S&TR��Չ��ɨEY�v���� 2jV��UP��G������� F:`��Oa�f�N��;�B�>x����t6����� �3~$�*�D�jwHR�̤�R7��,�p��vͪ��zGI�����a��T��QQb��D�3�P���l�n%��W׺���~fZ:y�L�����=���wyA��t���PP�1�X�An���Jot%̇	���kk�H��l��,((�������5����|�T�F$�{t%�f�b�q��f%�go�%Cy�9�@@i+$*�ƨa6V�}��/�X���W}7��ۢ;��&��,�U��Jf���)�yB`���K�:C��>Ch�0�V<����h��:�3���h���(WO����W�̀�����]=��.�e��&Һ�t�$a��ۚ�-�Gi֎_;�!����.-�Tc/�cO��z�X�#���C��/�OD�����p�΀m���V��+ϩ��ɅIc�?�1❵P*��p�� �X�P�L%HTDhO��ӠmGtZ^����v1�L��a/�Հ��*�\��39��"��A���Xx�#�����Жd����	���!a��q_6���}L� ?�v����>���N�P�iٮ0{8�&�4�/�����"�t�f�G;5/��) ���GM��Ѿ4R7�ܟ�y����[���E�p�=hb2��2d[���D߆�����9��5������M�jr��H]w	��U�D�i����V�HAk͍bJ��o�J�s]�k�G��S2���Ʉ�$�YU�"���`£�5ĊR�s���o�ٰZ��fT�?z�yP�7����������[G��Y��*�[:Џ�0���O�w�ym�]�Q�4y�sJD[��9�@��û�^��gE�����Ux� �e��<���"動#̌C4H��# �	0"�	�B����h�ΣrX,nV)kyCڅىa>�����7s+���f�jz~s��"�=�w~ʯ���3GVQ���vڀ:J��/BU����=�M{�+.� �bɔ(�a��M�y�)y	
-%裥�g�փN{A�&�=�iZ@7��o���$�7�(H#�� #����F�]�Vt�(��.Y�FE?fШ����of.t_:��^Q-*`�v��֮��n�rX��L�_��Z}��wfj�����cH־���;�2��Mm�L%�m���M_H�{k�0a��ML��a��-�`v�q{�m�P���!�4dl{+Û��Q�Ř`��M-5�M�m_����SJ�������m�����̻T��{m��@�F���@�CFr^�ْ�'���?�cI$�,�K�n(�v��n�Ѡ2�ݨ�@��z*��%��/�Sn�l>���ue�K�%G����_7ץm����vY�jV�L"�
�]�҅74Ϭ����Az�t'��"v�o�]a��/�L\o^�<we�#Ba�]�`x��Q���
�B����HX%��ͣ��%�:C����pL�Ғl�O���1�ua��ђ�s�0\;0������B���� ��"7+�@:l+$����r��x%9jӃ�7��ݡr3��-7l�	��E��iկf�hԊ�4~��Y�E�-Bٞ��L��a��7�ր,Ղ@m�Bh{���W�=�#cT�ǚ��v"&�&o�P���� ��q4���X�W��B����W�D�W�Q9���R8�m���DF��ݒ�쓈�Ļ��`qy��	���*X-�7��z�W���擯D�'��ng`b�t�G;/7^I��`�m�gVJ���X��\��Sb�����V�a���N��I�;Af:�]#F�-L�"�%8ؒA:y��m4��'���t:� "�t�o��vv�=���-Ms��t�/�qO�6���'�,�0��E�>]��S��K��yv�¯�qec�w�-��)ҕ��+����mtj�m�_RHw�Fb��uR���6\����c #�	ا�{��_�q�dP1`�$�r��!��Վd%\���U]�[/���l�F)L��ًO����D���B8h��_��eA�<�O��m�hؿ�/��	7�;�׹k�Y}f�Z�T����=���Fצ�͈�JƟP��^��`����cŗ���0��l��@�#/(:	�Dh� Ӂ.@F�:Jj��> 4ɕ��u���\,����u�Y}���ί|~l�O(q�ا�Cy^�p(s��NG��W͏������e�a9��}��,Vv���W���Y� �ڗ�/c�R�>��0J��	�C)ila�]��8���ƻ�2��M�T~+�`@�_��b�)0G ?��Yz]fb.�<�&B�ԖB�L6خ���R2�3�}N�J1"���M��Lq(-�y���"���t;K�6]f���]1�h/CJ��B�E��� ��:�H/�2m�ԯG������%�o�Y����\ ..ķNVaX�?9)@]�������ӝ�ہS��� &v��Qˈ:험��R�~���A~�66����w��~$�V�i��q��)�����H�C�(�/I������%�� �>gB~�;I�z������m�ȯ)��/��C'(m�	/�>X �`�(��s	�$K)����=�z�%�c�M���A��Gq��HY<�qH:d���� t�6�g����hh�]�z�EO��s�S�2(-�(�Y��-	���f���0�%����f�����-a�,z����_��y3��Li��Ui�,�NA��/����؟6wf�o?��slm���鮟J3�j�9Mw5��&���꿶���.SF�y����PRճ�62�?�+ ��f߶A�![�Nd�w`�����-~����Zm	�-���2��$_���8�1)$����0���:V��>E�m���fu�f�6�1&zS�;$����a*�*�sw�����t/u7�=�ꭳ`�eƼ�~Aї#7y�h�~�;{&>�\(I�^gf4�5hD�۞�$D��~0��*�`��$/�JZ�������BD�.�-�R,/3��=:W_�Jf�;e?�6G�C��z���*�k��:oK�1��S=KzN�Ӵ�cڠ��[���n��;��oٕ�Š��ܸ�����Ǆ�B֤ڤ��Gq��K�J���&���d�\/h	��b[~��_���Vwfy��6p�:����C]���1�"�s[H�_�?��nv��8�p���3r��&8o� �-'(z�1���eJ]�˰*�����M�nh�#rTk� �b�9��j�2-^�����K������m'Q;䇻Yq+���\tl�my$���xٗ+֤Kf]t]0&oex��~�6�F����淋���}�y12x�CҴ�������M��&�@����z��	g�b��?/_���t�ai�'ۄlzh�}����%�&&���ڀx���Ǥś�J/l�QL�a+��¸�A1V�9e�X���4�E2֛R�B��6�C���}u\:�@�<�A�O�U�s��K�Sz��b��ee��:Lm�tz9�uH�4����1@��e�Z7��n�r	�ocZ����ySH�L��j�Mv��8�M���ќ�.4v��$;�ub�����͉?mN�2���^��tԗP����q,�UN��Y&�U�Dt�m����`�����\| � lPQ0O�ˆ���l<��[c���	[f�̧���=E�x�)7bAob�A�����
���p�0(��F9u"A��FJ�0�:��D"p���sd����Sc��v�#y�
�%'�+�Te�eo�M��Nh9Y���M��k�X�c�P�����z��r����#^�?���k��v��?����/;��`3I���v�%YΉ���z��f3/za�w��k�L>�������Q�b9tYg.���h]ZX��)��%hk"�nBԝ����S���P�~&͗�c_m#��JN1���Q�D�O�^$��|W�νSt�$f�}F��0C<1��4��W���D��F��-���	��ʥ�Q�DUo�R�AŔ�,�s�Lo�2���/���J�f��	�h'�����sp�'2���
��T��E�l/�2�7RM�C=A5��ߵ`,�=�y?�/TF��"�w��s�L.8\�"g�P����t�Ǣ�\1�eHK�����"�G�%
�e��L㓃K��:Y��(�GF}��>SѸo������o��q�(���5g�
/�lC�����?ok-���r����G���A��8	L2�ȝ��cmUEFJb��mS�a��*"��C�=1]�;C�~�]�����Ƽ�����..�E�l�0�f�����^`�()/8�2q���
x��v?��Z3�ٰB��4]8��Lw �G� �+jf�y{Qzم��f4KЂ�ܵ�8
)2��=;&�j[湒�Oܜ.ܑ{�s"���F������D�RSkm�J6J�2�8�+������ְ���$�sW�����_ȗ�wk'��z�C�  ��t�^�m�~h�m�M�QBU��K����� �\s�ⁱ��.����[��_��;xFDl�s�z����D�+��&�l�Gp\iD�o�
(��'��pym�\����V´���IH[�?�PM�I��+m�-{v;jJ��FG�*��32;��ۺ@������ܐ�?�������Ė��<h�V1�.
)����5)-���W�w+)cLZ�� X��V��8-�/9���ә�i.q?����#�����r�2�}��g^Q�i��6R��
��i:��̍p����u7�1��M���FU�-{:�Δ!Ā���j�@�,����! �}�ad�!s1[y��+D`GQ���)ezHa�k@�A�{ѓ�A85�d`ߗq�K}sߖ���6��]�u�gz��}V~���i�a�(wH����2<��N���';���fJi�9<���(T�M�D�ߏ7��T؃&���P�B ��:-��ko��.��v�=�%5�|�+X�����/�߄)��;P	����kDA�d8�(�M9��-(���W5��Vs���㸇�PP�}qH��u#(z���p��,�#����h�K�f�H��ZI����:|}�?L��g�����b}II�/�&� ���-t�)�W�01��k����W�2;��K���V�*<F�JN�n����Y�HT�e+M)8x�s��`:������hZ�@
�_��%'.*�i�t���r��׶�W�[(�v��dV�W�ӊ�Y�ʺV&n�)fӏ�`���^���\'�K����a',�f��&�he@X����-ߎ��n!��+�O���|���@� 	��61��6l�����(>QI`����&V�*��cgq�G���m8R �/hZ>
����qjp���b٩�x OXp�(�)	�ҕa�������?��s�� ���Ss���ɶ�[��{���t�5)"��#�A�Ƨ�q��`�W!v�Ψ:��1uO}��K�0����%F0~p+����sY����r�l�%xP4AfY��L8��#V<�z�+������'B�/́�����h������ꤤ�}� �x*��'��ޒ@tRa	��@�*�
L	�I��l1�y�ﺛp�b���$s�T������й�;� xf�6��+ݷ�ǶƂs�Nx��lr�r�UpΝ-�Юw|c�LH���?7�.������"��t�4RB��mn?p��!8�̂�׳Б�~n?�U\3��;c�>���t"�-Yٮ}�&ڨ\g����q\�o�}b�-4PN�,p��M�upw��Aٿ��kƀ�ں��U�k�y�ؤ&���`�f'+����o�ioc$;�K�G�JJ fǬ�׽�t��)����U�ԕ��9�k������(}����a��;����:E� �"�� :Ctݯ���P~��I�{N���e��[D�'�"Ć"V�^��Pg�*�hn���j��zDF״��޴�5n����I�;a4�s��?l*D]۲(�b�E�ce�nYގ�-6%1&�E�1�C�^�ݒ�h��`���L
nMd��W��+�C����(NT�$X�����`������e�����)
�2d���9�vZ�$�385j�wE�l
���I{Z����F\�/ԛv%'L�o���@�i1��Ԟ���O4��G��#��� ;���J��#���	f��m)x_%�⸹��S��3`�����:�r�镕�ŀN�(o^h|����ĳQt�.�=F�����g��W�#p�����fãs�i�c+�R41�q@ġ�`��S�Kw��F Ԫ� �����^`�&���=3c�ᦴ��%Au����j��S�������-��I�<~p�����5̏˦N@`eU�}j���e��>��`g�M�j� ^��p����XB̢ [��2��7t�˻��+�{tش��N���'�沵SƵ�����O�'U��߿��ذ^�l��2[� b�G�_��.���|����}�C�1R�"�}��q�D���8G���(��"����Sф��a>ޝp�&����eװ ���ڑ�5�_�v뱫/TG�5���#������UU&�}��vk��~X$Gq
?4ۂ{P5~�I+��?���8"4Mڧg՝
S4�օ���(�M,_�v����,��"T�-�ݓe��vN�.|�dZ��H�����`|�м��U����IrqN��(Ѩ�Ew9h���V)iܙKN���ԑX%��T����1�z}��4��}2�?cB�F̢j�(%�u�^qS%���`7�����(��%e:���=
���VO˅�M����Z�!3���?�ïB{�x�.JE$#���1�3W�#TL��<=��))ax���qz)�o!��S�b���Xn�l�4�Si�nۄ�����h�k�Xifl�5_�F���%ob�������$W]M|{�p{�Z`�\�L�Nb[��@���#�y�tuBh6e5�I� Ad�?����2��R��.�ڢC�JcV��F]����zyVGc������/n~�T�!��#p$��{r���	�j�ߺF�F�8������^X<<�n��*�d(>5�!�@zs�;�Q*��=v�e���0;�tEF���W��-��^sD�;��w,�mO��D�Jσ���\��-H�"L�J�Ⱥ��$L*�����*��d�&!��M�!�a� a���I�>MK���vT[���07ڑ!c̊{c��&V=J�t���z��<�!2o���d�E�ܡ�i����ן~�ȥV�3[!�x�����/q�y|���"����)F-8.��[+!��
(�����!���G�y��g���"F�v�)�P���_G耩a�Ny�T���v5'�,55��� K���t����t�k�N�K1���#��K�e����W��N� V�/��P�o�كӢ����7��D����Vv�w`�vq��#F��8u�3�jUԂp���ٷ��`�r+�������� ]p����f:Wy5�f��sm��Y�$tj��>�w&�����OĴ������β�	�y�%δ8�Xc����Չ��k^�@T>:��.۩��#*J�컖�{�麩3BUQ��=�ҋ�+�ai��������cI6e_�i�A6K��,�2z�G�
ar��v��1���~yp�w0���*F��P�.�f���x�a���"�	��b7db�2y+�l�hP^'ۓ���#")���[-d���<3�Ĕ@��}���ʜ��'_3n�V�^a�V|��f��]"�l"=��I���h�)���B��i��`>�n��ы��8�k4��˶C�k1��-<Loߛ��2i�,�O� ��o�YJ�SR������zt�`Z��W�H�	�
rܑ��qֻ ��ʆO������JK���,���qüS��s�v]ZFG<-���6q�!���Js���
��]qy^��Xf����E��{U^��G&EqӠl�a6��u3 ?�}���r�2U�D����4��uf�s�;K�M�'�i�՛/��L�ӈ&0�m�ޗ@�U?����ғ�xR���
���S�/�ynBxmE��{��Up�8{.d�\��9x��Y/j<�_ޛ�ƶ�?���� d�#:�����eo�ٴ#�(-"T� �@�[$9��T]~�F����NMW�[s�LM4%�p�)ŷN���ө��b�-]�r����ܲy.�\Ŋ|���ư	�D!�S��pW\|��ٹY�[ǂ�!�a���j��u��n��-�-A4�6�ފz%4`Ɋ1��	[|&- x��2Q�ø��WE�C��a#�����l��������E-0<z�xio�V��	��=S��d�}�>���;C��0�u�̀��sC�u�AcP�L-��e�M��#7k!�Kt��2�_��T���a��$弲N8��� 1r&Ʌr�G9!ɦl����Dx2Εa�%�맙�y�&��1���H�R�po�Z�J��Nh9a�-���&Q�0(��XJm�g��z���`��"�`܅=���LS��'����~���-��L���(i!�K�s1�p��d��/e�� =�Z���"�z�z�1�b�+����#�w� ȵc��PƒWjr�}8~���8���K���X�v-�<dL����#��pY -I���Z�&�0�׮^��~�:0Ѱ��LA8���%�Qo�)>�g�:^�Y�Q�Q&=�橪*
S�J��}EP��	jʑ�f��E��iM�0_��IfwsY6�wh�������i������Os�=�	s����?u;e0��QI�Ʊƀ�|:�R��`�X,C�U���5���}n�/ƍ|T�}Q����v,ɹ�rx�A�9����̤	4�<Z2*$ʲ�	"w�b��]�0@ ����H�T�ག;K>=�Ya����X�TxM9�Gqڨ'�-���*��X��w�)�:�#\1ܑ|��qr+��n60��v^M�]c�lK����u�d(W��r�q`t���lb��:и5]��x�3������?����A����`��/I[Z!Y1�,x�L��7�ϧ{���0&�@w7H�w�����Y�X�{�}�Cc�0Wа��`�V��!ߵ����Չ\�R�3��cqa���j��w����y���ZDs�vf)�ÿ�{	:��<�A=��|��'�(�4؏��E {8֤�k�z�l<�����{>��%M�`˻>I~7�g�Xq�Y�h�}��ٻ�p��/�!�:�^�J�l�[�^�� �������#攃�/ϳE��}�����>��Y<���]��{��nnX�,���d��(v���Kb�s#��Un�W	��Q�g&-��i�= ݽ�J`J�%T$�l�UԪ����PA#�h�:��VZ��D��� ����Nd�="�z�l��,��`���`�Xy�#�Y����1�C)�$MC�z@��s�J���9z]�~A�Xf;1 A�$���k+�
��3!(�ݫQ�ϋ�PB�uP`�6"(�o�g���e	�`�i�|0��fϡ��dgO�%��cZ�,m!�ď���Bġ&[J�9�%:��[́�� z�W�lg�K��	��F���a,�4u�&����C�)C�6r��@�nm�/�j�%p�g/���H���¬`�q�?U8Ô��{�y��$iV�y����i%^E������@ȕ��n��H���� }S`��I/����:�ﮣR�ز��]�9�/�S*u�ޡlS)��ϗ�"�\�\�`u�|�!փ|�TA�=����ۍ��1��9R{�륊Ѵ8Y̛��<)9LP��q������i �0��$ e�G=?�V	$�����1=d��K���~q Ԁ�ȴ'PV�/��ex�[��/��Z��Z�����U���T�)�L���2+��Fj}7��Q���.�߹e�"�e�a�A�M�f�+��G��o)��#n������o�-���7�"�>� �I�p� &B�93�XF�3}�ubI��� C%�����&b��d�TDfAy���U)��-���q&X7��q3��w�:[����3�
�Hm���c�e"W�9�F"�>�..@M*�D��G1����ca�x��s�R���L"�q�Ӷ��`	B�@���
�Q�'����I�>��
�J=۴�����/c:�;h�*�o��݂�3.j���1��g
����C����%ΓW�L�EDf�Z({�ԑ��_{QY/s`��5���P�MZ�}E��T���V���fDQk�JYA�Z+�����/v�w%q�?Ǔ�t4b%W�{�,�d�W.Ⱥ�Ӹ���v�(N*s��m�otB~8 95�fz ̬Д��W|k5�@ (�Uh�x��	�q�pH!�M�w���)���*��E� Asv�8�!��Ǔ��t�Eg�5m��`�������O��t�WcN�\�e��R��1v�y�5z��"q�mL|���ml�=���~�6Ó���\y}�J��*�Ƈae?���A���A9Jؙwy��}E�ؙ��gZ��J4�^-��6ҋc��Z�nF�S9�d2Cc^�0�`S�FX)���3%�����tv�iQ�"��u���h��;��F�<�_��V����r=i4�Û���jtT��JCS	�C�77G3Zk��_hH�$ǅKl!�7j�����ן"u�yD`d�(��r���6�]�e�I�edU��
��T����$�php�q=4�[���ޭ<��g��+�Z�N���&7��_�ʨ+J����6z�_{C����nus�X9(��W&��`���^q�.4���`�qE4�+Ⱥ&-jeD���/i�P����/ �F�&!�>�6��_�:��J�{��֘�m�:چuޱ�KS�>�+)�ϟ��pt�C��U�H�A��̯t�1�W%������ۼ6k>W�L�f��Qz�h!��a�ΐ�[�$y�oC�~E<��i L��-��X��lnS�n��XB������ņ[t�m3V+zwb�wx�Q��p ?xߪn+���Gvr�+fԟ\?��}F�F���Jn+ lj�Jzn���=	�:��'S.�U�կ�
�b��`��@�_@�\��c�`�,Z������n�MxJ�5<�]q���#�'f����#�ܵM���]��E�١�t�+��
�|/�$t�8Y�ˇ������!��#�q���*�]y���V*#;�'�a�&	�i���S����J�`<{+�rЙٓ���;�v���w����@Q��{��q�J�h]�?��I��R�祿��/�grs5wn�$u���;&A*�JA�<��{���8-b�(���>k0'��\�%��A@��ڭ;��Y|Ag�mp:�U��3��X�� .RM?���B���mML�]�c�ԴA|3>��({e�]O��H��6!K&�5=3�j�d�%��k�ِ�R�R�3��сCG�c1��j��\�A�ep��|����/���#�y������3d$fh /d�!�	�ÊD�4r�g���{����C���8��W�ʲ[�f�nu�&|�pĭ�lH�S����W�h�f�;�˯�袟�-��p�����8lmMP�l؊�Y�%�,�I�8�@�;q�{���u�K�E�q?���v�ţ"��*?�ni�k"\+���Z������9���6��c"���2eIu6N\�
�b�'���p9&��E
_��{kg~�=>����C��(�泽�0
Xm��λ��{����x9��*�Y��q��*� 5��je�,��K�ݙ]zŃ�nX���Z���~���$�.��:qd���1��)��-����Z/V�'K
툰��1��^8��:-���֠�_IL�<%��V{�il�y��+��(xi^1Y�)���dv-_$PƹԀ��̰��o���k��h<��n	F*r����1��ψ�|����%���H^y���T+�)���\z�F�܂1)ܵ�E��ޥ�x��a��� �Ɖ<�x�S��ۈN�+N�v�Kq��%Rh�C˻0vL�����9�]���e�pe�B"g��T�)=��_U���)l"�Yˎ��Y�)��y�3@K��`�#���݇F�E��G�+�o�OlUK�x/w��	U�ၚ��6k@�8�;˗�\5���� *ܺm�myzt���6�z���X�[�@���m��tNGg�t�^ �i�|a!�A<>e	M!"""I��㢃胿���U����������
J��mG��XCiR���JX�{��(VKB1?3R��
�T/�<1�������&
OZI@
�����U�n�B�cZ:���qv}*�W�#�}�D�+�u'/
ܤ�CtPm�&0�^O�עs�~C%���L����d�Zb�وI�����Nc=s�'%Cb`��y^�@èSUU^�՚~L}����숈�p�%O-C��}�d�JꝐ��8r5CR����[뮃�.g�pW}� ������
���f����=����f�y���\6�⎢�OM�p�����Gc����Pd�a�4".dvT-T֛"u��U���p,�$Dy�ZN�yF�ФV�N=�16��U�a���d�kr�Ɏ,`�BJpn�<�/q�
��`�����y�r� �r��}�$��VW�:[Wt8���g@�8r 43�B+̠n��[����Zz�,�8��SG���3��ú�N�K��*�5���j+�Y�t�n$R��~�Z~�J<��t�ɚ,�^x�D�.}@w���d?g�Yr �r_;��M� x����fL�GC��dl�P"���f��X/�:a�d�#a�k���\f"��Z�U@Nί2���̋|{h\N&<͞�����r�8�DT �/�s��1:型�h2�G\	��ie�˗Z�ӣ,��u��^R��w�7�D3���:ߊ�3鹜��� �:f����賋�-
�'�
���{g�Ƭ�ġq*��IH��T��Y�<-�0	�3㡆2�Ӿ�Z#���??����BM�4l�����v(�&
Q��F`��t{���Jr!���HR�Sy~��ۤ��0�.<G�Z��<$���LL�:�P.T˿	�ϕ�bqi]���S+�~���$�?/��!&�'>n�с����gJy�$�6�w�[$����8��Ќ�s���T���O>��u:����a6Y?xBD���FJ���g��jb�> ���]f��GD��[+�G�����%�@}:�At�-=d���^~���_*3n��xn��|��>f���S(&�~�[�sل�d��� ����b�V�SR '��)���D��=�J�?RRX�*�F�C�+��zHL�~�V3�{��'5e?��c���h�Z!�E���Wv? ��t��sr}`����j��ҫ*��a�T��$���E���8�?�����X����[����a>4��
oN�PA}Ԏe=b=���%x-���4V[��-k�R�A1�Z��-��J�F�5�O��1�	e�ȴ�2/�Cj�4��D��g�n���4���=kH�F���������4rd8���PW�%`E�F�jW� �I��Š�!#a�IM�2�{k�%�������F_rڲ�������2��';"$�r�ށU/�Є:��I�9��eY{�w�rX��K�R��}� ��KSM>�Lh�k��,�!�����>:������_�ɨ)���Q.�}\��s{�IE9eԞH��V��DzL�r�_}�\�Yȱ��'���և�s;J�����laQT��3�F�q�@������r��pOg�M�T/7-��PH�*b�UU�8�;�(��1$�]�B����O������7F�!4k�C�x���י�Mg<o�K�~�6�5� ���&�����ea0`�g6E}�`�����s������Io����㷵}���O�_�_�� )G�ᵇNo�_�I�1�����m>�P��H��٭!`|����l��7�<y���Ŧ�Ww�%p��4p�Ty���2X(H�i�6ku1�F/��S�ݾ�kn�Ȧ�7�D�{-�nhp�d����R�#��˩7��i���d�=�E�R"���S�;�h�Ĳ��Ȱ5K�2��m���z��M�T&L74\����@��������_%���U2O���/�;V�i�8NCe��ˈ1
x@�/m�U�S-ߟ"rg"U�uw�z͎@t�38�/�pr�E;���e�YM�O���N�Րe�Ȍ��Nn.d$���}���Y��S� gi�o`���͛�b���-�Ym
�<���$���7�@�Z')v<�_�Jl��D�)��[d�	ʴ{��F���fh��]�kf����>ʶ�v�xn�KK�.7���%`F��m|�ٔD��Y:>��7F|���w֘��=]zZ���9�{U�n���D[�ǆ�Ƣ�29ȡ�}'�p��r�N�(Q��8[b���<�Ck�^�����
; ������Z�D��G��.}�� }t��Z_2q����Dq�����"��o�rj��"��L#*߫��C����X[�?Ƌ<a��A�3��������(�j�b�z�gc��{�t@4���'N�d3��az���	����e��3�����
ڌ~YULV��i�@3��}�!�6���b��a�@�����`U���HM~KXl��1��FxeV��ɛߗ����`�~����喀���#D���ێ������x0�ః��ttP�h�jM����i�4Ѽ=��������ש��؝����LĨ�&�	��T*Qk�>v_cD�An�-X�׌�.��Ӌ7���o0�q�B��n�ut���*�{g��*D �W?���q�D�gq�'21B#Kc!Y�7��7�n�cB�����ͭ��S2