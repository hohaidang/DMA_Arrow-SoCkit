��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z�����4��������8xT�(�h���/�<�F^[��V<v�Lz�=q{���ˁS�=Y��y�
��+J7�‿��(��ߑ��gƄ���'�j����/����Ǟ�H� �a�C��O�m���I�_���"kI�Sο�!t�Lp��x�7)���2y�����d� 9��Q��Ԩ(Gl�G�-�z��?#:�?��>��R:`: ���X���g���&�8��0��	��ӈ�d�ҎQ9�2��=�J�=��ވ�
EHC��M��jQ�����7[<jQ�AM��S�r;�ZP{2�*
�k����ז�=��'�����kBl]�lnyg�x7|k�f��s
�%arϸSX"U�-Q���� �?���*|0��|�;f3SG��{�c����L������[� ����ek�����H<�EϪy�3�ǹ'k	A�wE����k�jxxZ
�)bC1s����t��vM��������n���P�L�7a@�mMixb�F��X7Hr��-!O�#t�_vy�ɦAƖ-^*�Jp��G�\@n��24��ga��&DX��~�{�W�O���(�Op����%�<�#�W�rp������r�w��P�j�0+z�I�&����!�j'HM��f��F4cqW�3g�����W��{J*fB%�>+F"�Zd�=����E���5���U�H�$�H���4���ǵ��X�tW���	�����hCMݷc�ֳ�V�*���Ej&CT�U�3*��M�d{�aTf�u���8E&E�s�Ϡ���2�$��x����N���7�:��S]��c�b��#��93�~������s��y�N�
�	�r&����
������#�C�nl,}�7�Kq��� �CO����I;t�g���Y<_��C�����b]D������W�iC�=e���9j�洏w_3R1�>lCt汳G��|�n����W�Q
��}x���̦6OfK���;�X౾��o���,>.Ė��uw�
e8k���6����'��t5,c��%Mb%0�C��3��!���6�ܪY˵�#��:��+Z�[�c�7�K��Ţ�	���L֚�ۏ^=B�ׄ�|�+7A_���"�H�\A�r*)>����!���9r
%�"�W;ߠ�FOkt0u2A��<�1�uFh���
f��.�:`ODXS↬:�������Z��)�խ�5��|�us(I�b���H�6��G�)[�nC�$�����8��l*t���&u�!�լٳP�y_D�q���� *���4:C�����XOn�i��'z�<�Z��&L���m���%���7�:.F\Gq�W_d�<�޲�?�eۢ�CḕC\(�<7 ?����*���H����K���DY䯕�&�O�U���lf������d3�6�2aQS�S�l�`���S#*��j�ɢ��3)�\�n@D<�pU�P�i�x���G&i����[ޙ����|#4��/���u��+~�	�ݭ��z�{<��ü���`7�O��x���D5�o�9}݂)~ �5�2�N ���2�I�ZI+[|\���.h�T�q����x ~<�B��g���D���7S��z#�P_M�f%��Ű5nr}O���ֿ��P7�����p���
��("kQ�	�>B�rr,�]�A�X=�^93��k�Q�Hb̚�A7y��B��ݵ�����&�.F��ˬ��?�,�Q�Wi�63�X_(�s�[D�qi(m0�ʠݢ��8L�oKous��
��rY �$�Hi�E��{� ����QL�6�3�lU�҉
�]�dASZ(D������t}��T^j�
Ue�rvq9h�<����t�j�!h�5��짮E���϶�vj�2�m�r�"�XS�ځ����_o�;ne4�-D����S?
����m
�	5M���h3��+W��X��N����=z����i���h��1)8*%R,M_�MQ�:pC�a��ʉ�^��aj�O�n��G�7oy{|�jM1���5��P����_"ғ�DEՌ�
 �DW�)
�ZE���9)�.���k[w;$�����$*)�-i��,�u?z�ne�\slh�Y�*��h�!��b�67-�:]��&�`�v�M�c��r�.!8�������[�F���d�ʞR����E��Cg��L⨅0�#zIB�_:���c�V�J��v�,��$���L�S^~^z�-bb�2՘cY3���T��A�ϻ����O>\RY�pw���1�����#5C�Ybz��2�0�-x��8�~=mERP2)FV���g0�-7-_�V�es�S9�68&N�Ҍ���Aݯ�ʼ+�0SD�e��O"��⏏��L'yR"(�w�h�-D��=x���@v��x�0�bW���3����p��W='?���z��WfIlQ�k�T"d�l�K��w�k�3�Kp�� ��Q*�[�
ѻ�51��Ks�4s�pB5JC���ș�M�e����#�Y��T���� ���"�۩��)X�0cyn���*q�&��f�� h�10��;P�cEu�
Ƒ��2�*�YVG>�k��~4���\�Ɗ�{�V/~68#{���B�xB��!��ˤVd��"�H"�%Úe�v�h+�犐�/�8�}�q�za�(�k��G�l	�!�9@��X�ь� ]�dx��9+Yl�'%��5��%�zi4�u�{�2}��w�d������l�%R%���#<�!�M�~�+�A�r��G>^4�4��8$�3zh;]��x2�H"(e#�>��.�H��ٱŨB��TuEd�����q�Njɝ)�Sʝ���ޖ�4j�
�-�e� Q&�*���X�	�K�����8ln�*v|�3?��b��u��)";zl�e�^�/K����%��0��Q��f�](B��p2�	�q��(�����m��&olo��d���ӭ҂�<�NH��m�����]r�[��kw�zríS�_�	 ON^u�`��ؕY�X�4I(�Za�+�C���������׶@�0��Q����Gwu~dpABy��}PX]�����SH�R����=(0ؙx��3���t��֦�dAA�h/*�\o��g-5� ~��/���/�����7e���6���_y�)�[M�e�,M�rFAL�iF b�+\'?UI`&�2��5�
�\��0>�m,�2�|��>;�T�8����;Em.]�D����������~�&��X}d�D�9������^�ku�_+����6����wg���6uOP��L�|OP��'�t}'���E� �*GPc��.�_5Ą*�UFzLS�5SgSu�ߗ�\��c�ϟ�k�w��L!V?��j'm�W�D��l]�h��aS�I\�Th͎t-����?�de�bʝD��۱��]'7�x9�\]ډ���>{!���N�Ɂ�E��W�	�S���v� �������op���	�~
������9v<�dv-������`c�Ȍ�g�Z���!���k�KH��W��v�k7��@�O��d-��;r���S`��%�U�p�=�O�$d��3��iXk	�[�����aE��MO<!�%t~p�9%Ӝ��ȞH�<��xE�%�-�<�}oǳ�@_J�Dr�i����oy	�u�=3;�ͭ�W�R��Xr��ZU���6:�겦(Ψ�����t�+|B�9n�0�$��1�n�S	�  a[0��q��Ĕ��=�k��5}Ze��ije���Ӟ���D�s�M�)��{"q)�2��aN�P��Cy�$�j���ё)Ϟ�>]�>2�.���H�{�{����Vr��[��K����{.�0�-ə��f#6E�(��x݃Lj��vJ��=������+{�zx&bU)C���ލi>/��]܄�=�Z��s��n���� �$���R���JO�N6.�3bL��5�	�<򏐚�YZ�@�������?� &n҈E�J�Rv��Ғ�ś_�-�J�e�}����P߼��G�z���S�y�EE�L~��\}���UvX�"$èX!I��<�HaV鰂�+��B(w�I*]���"H �]˫�T�L�7儦醝�z}/1A�t�$(֬�a�@.��kyr�l5�h�3�1+$r��ә�V��� �"$ƽ�$��՘�Ӏ�t����^81+�r����S��x�R��^��������م����;��W�=H�=uv=t��?�]��L������4��D��T��7�����J�^q��,D�	O��Z�.�<�	�%���ʡ�N\by�#w����澭��Α�3Ad�JB�jJ��V�j�Z�4ϩI�:kH��,�����9ů��;k���k{g,�����z�w3�N�Ǡ5 �4��o��Lw}�$�c���ۊl/mx"Y�,Ĉ�ō6�z���SB0�;�Rn�b��~INÖ
���x������uE�5����	"z��Z�~z��1�W�6w�+ǗU	�ق��GY�^S�] ~D�|��Oq���c2{l���rRsu�.=4��I�܀��)����|��D�p��� W������� D�`��t�Nϭ�����tYN07�
��3ZO�����O8�8�g�@Zy#�m/C��P��9y/uw�V����Q��v�� �chp���>o���3��CH �APpϠ(�h'0 �� �eC�i*���D�}ئZ岶 �Z���:!:��r��^A���h.,�:Z�?�җ"��#9H:��M��]�������_u�C�F�ޓ�J��~��o���+ڈ2�b�{#�"���]Х����~]�/��̷Vw���18iY͸p�4���,뭟�����$��@+��`4��B)�>�\& �ݥ�0���Q�ԧ��x9E��ɺqU����c=�ڭK����'P�-���awȷ���lx��0��fT����P0(�����L��%��?- 5,�爴�\���\�����d��!�(,c�ͽROC��nj��������J%�\������m��a2wT�Qݧ17C���I�Ss1��S�@���֓�E��PJ�0ڌ������5?�d*��\MZ��8U�3/�� ǂ�z�~&�����L�|ܶ���ܝ˚"�2����g���[�iZCr�zp�|VtpH��N��u�ޭ��9l�w��n,���#%�n7�	�i@@)��������Z���x���j�"&sG�H�V�6�^�E���V \4���e����k��'��a9O%���&�������/�P��$�r����������D5�T�����>+T`� O�A,	V:
�~.G�M̾m1��ҙ}7t��hB�&�paq���܁3�`����a
@s`XH"�)9�.�sכ��_\ب���"��.f���7�_~��r�'�L�lK��R����ԒW��� z)���U�jZ����d�m���z(_ЊR5}����9��U~w,6䛋�ye��}>�V4�<Fl��^gm��D��y?�#�}��G�͖%%ι��,-�U�fq�b�����w,k&�,��$����v��dg�"�D�;Z3�B��4F��K�Q�͟Q�oq�B���ְ;w�l�0ֿ`}+���R8�dU���J��pڱ·�=�<nV�?6�)�.�{|��2u�g�n���8Ю��l�(�h[�碩�-wWP�v�����T���o�]�Q�'
����_52u���\޸֛t\o�b._����K��cjeb:/�M ���%�����}�`�;{ ��n�^�BdB�l��\�u靦}O�bh�"����/��Z�߅���u�FN0�OS�8�4���w���SŌcI�D� ���<�!WK�o1⍐0:��;(Y��(�{�.\v#Cc���P�֎���x�n�H�d�����8��er]]��*(�vIt�/��fV��ؽ���:;i q�(��%��A�>�W+6.�h������������!�Zd4:c}fjz%��F�G
PI�I��Ҁ�pơ�Y�Lnǁ���>�_˙�2P�;���߈���ۊ��N���������¯JZ�&��Dҫώ'��
'4q���Fj8�F�6�!K�|V�R6&�7�6�VY){rua��4�J���Fj�f�j`a	<'aƀrq�u3���h��3��:t���~��o�E.�i�*��i�y�؉�#�mC `��S����a�M���ek���b�Ft�IF�<��N2��OJ��S��e.lr������g�(�7`��Q��k��H>
/FP;o?=$rA�Uq��1��މN�uI�Ȍ%O&]��+|5k��o�iK�Q���{��F�(�| T��ı��D$�h�{x7��:!���5�1���ג��#uBbF;���+�cvB~z���?�\�g	
�7�R��{�	Peb_�Mp��"�8��_��nQ�%��Dg�Ӗ��z��~��⎘��u��Ip8;��]>�T�ភV�}��J
�䲤�agq��!�F����P-V��n��#���������nqCE�X�(f��C����	�)�_#&{\1��BpT��%�4�>��w&�^�"����� h�1�
�"�."���ꁩr����xe���.�x�b�����]
R�k�PpWN4���L��j�i�pXx���_׽�c�9<�0MvO8O2�%�萡 �܆1�(����Y���.Y�d�����ǟ�/�m��m��T��V͂P����5��������k6�FF��.M�ī�__�����t��WG����H�X�.��+%�4�9��tP�\�C�4ڃ���T��%��XiM7:�Һ%�Wy���#7����CI��0 �Q�p��0�,[�o�T
�Oα���Rg&
�� c���k��%�������7���!�C]-��
�w��9|	�����ßA�/pث������FD���1��A;��6|)"�n��+�-�O�=ްɴߙ�n�6������=5����/,o����"xmǿWQ��Ư�]���v�8�����X�*�17Ŕ��`�ǁ�AP�z�?��&��5�:ї����$΀��~6	��/:����o�������������һ���T�B��lN�*�'����K�.h�n-n��=��f�VagO���a==�tt��.��ϛbd���*��=W���L��X�����s�o�)㒌|d��܆|�\��ڐ*���K��G����1S���
��᳑����Ɂ����H�����=��Z���P�r�|W�LL��9|��43�A~G9_/��)L�yGTPså*&�8�e�~���DI6�}��؋�v�&_7(}(�K+��!�&"���NI3�����D���T�H�������ŉf���it��uM�~_��ᆜց#r�����c����I�Bk3���(W�,aq��1|ĽH�����k���bqbα3�2Yq@���=Oۑ������e0�ڍ8�
���F�!�W�>��Kh6��1�g���d�w%e�Ŗ�1Z7��z5T��FT|�X��F��T��ŷ�H�n H�H��E��'��7i���`����?a��o:�1{���\������j�	/��C����#���:����Sx{{�<��/ת~?�F��_��裺J�ͮ���/K���p+*w�l���v� ����wp��B�l�!�a{o��I2Q��/M؂���a�4I���HB�n��4st��W�ʟ�9z��nDR)�,�%���j�D����e	DKx ����8��eXB'�tN0�����7�B>T	���o|��C��S�}4��m;���������[��@s� {V̽��Lg4�(c9�;_�)���s<\AJA$ec��HǦ$�S��B�00���E7%]�f�k��z���8��lI�T���U�'�����Nx�n�")�{�'��W�)�O �P�4���r6�Ȕ,��T��`�3�M�6V��v������(|r�����x�Z\i_֞�0�X�y܆뤼?Vը?��� �Ϧ5��y7"���I�1Zl�.Ɋ�|�c��	���1���uA��sv�K� E��I�"�$(����V:f�	���*�f##��&%N�Z�0����Ù��g�&�#�!0���1^�P:��d^b�X�}�<��<�r`1s�c
�&�Az��k�����MS��
 ^�jY��&��	'K#q1����!�k�h��z3C$�PR�988��U"����/�3_v�R��4���V[UIa��r�������r>��G��l���Z��u9^|'y�y�!�=�g%�|ᙣ�
/3l�(�o�(�ΰ�}�F
����ʆ�ZG�M�Q-�7���	����Q������ Eܴ�:��z���B�W%� ��j2����Ǥ=ot,�����5.��%����L��}�ʤ@��a㤞ä��R+���X&�c66~�de���lM�X�B��.ك
�2�v�h�3�u@�� ��S��с���L?�)�7�j�P_�ϫ_<��1�]1+ÿ�c�+H�ù7�5,���e麇��]�FNE��O��d߄F��x�����L)��@?,ғ��|$�l?d]_����AQB<��
__\�Tۤ���z�Ͼ�{�<�Ȏc�����c�[�rKd�M���1�8��b���]��L^,��=y�3������5�PaI�P-���W��N�|� ��L�7m��C)u@i{���v}eʼPՌ�JJ��r��j9t|/9�;u^�oleeaRmn�Vf��Ft��ɩ�pҰr��8�iB��2��=]j������e��Vt��d֞&P��=�'�_�9K���VS��/'ۘ;��iW6�W ��P}�nմ"�l�N 4B��K�ȴ��@<o�=2�p�8�E�	�^ ���r=�W2^pb	w�K��i�nw`���,�/Ú"2�M2�'��@��遌c@W�&>���xӤkx�SX��u`NS��ݾ}�a裋���̩�ym$&���Z�m�8i�.����<���������&�����31�P;rݰ�ݾTV�Q���+���f�en�wʉ�R1�p$�d9��7C�]8{a��f}ҿ��)�܇Ӊ�SFCZ�VS�����FνEG������"D.��A�dɤK0�&h�lM(T����[��F�Ǭ5��y}闞��t��cm��6�n��h�cs��[GӁm�<Mi'N%��������L*���^a]*`�g�I�c�K����H�O�NRL�s����H,�ڜ�a�S_�����AB�}{p@вnPU}?��&Q�ϛ�`�X�(�GKR�Jذ���'��R	G�̲�c.���V�Ʌ���6I·v��E���I �ö�|��u�Fۆ�]�;�$x,f��'�i�lh=ƪ�5޺��Au�m�`M�b$�;�y���u����I[�(��.���g�Gc�?��:��}<�*�d�Z'+��2;����`OA�>�}���˯o[��Sg������t_�B����7�6
��+e�@�<�`��A>]�wP9��Z�j,��䢟�.D�#�B�1�;���F2ȮdG���`�mht��y拾Y?����jrd��o�?˟3}Hx��<�����IW@��wg�2�.����&��#�O�I6���#E��v�R�
���?V<��M�� �|��ǡ+]�	;���o�E��h�8|��,{D]q�� �����/�r�r����5}�q��C�N ����� ���F$fbD:�'�-Hp�=�o�6���~�V��{�{��Y_"�!t�/�3�U��{�|8�tpA�+T�-����Z���d�E\u���C����;�h|�P�<j��?���S ��ԡ+��Y^2*�<D�j]>JԜ�u0ͤ'֛x���i�dΕ~s#�d��r3���"��3f�K�
k��L?��p1�c/CW��i]�4j���*�l@��/D���G�P&`��kyܰ�;{��-,�6}�:���m�����N�&2��Y�z�}[%��6��v�M#��Dk�N�w����<*�{����-ҷ��"�B�G�v'Et���"Oy����Lc�5��t���[�!v����@�+H;�a#"ɔf�Z޵�D��u p�N�A&�:M)�pB{0c��"���=���XM����J��:��5�=f�ov�Tu��uh`H]��=ZQr��T�/�F03w��T��e�c	���Z�J�����Yk�;�L�yi�%�ZZ�`���n$ŕZ_����F���+lP;�
��BSS�j���ڞm?�dR��2<aKQ�v,����d7�d�S��ڳo��>�i����;��D�+�߉�Q@�Vg�[��/��Hw&Y�y��d�)�+�%Y}O)Z�������)^*�9*�<��}���tz��pFPQ�4Jv�6�dѫ[{x�*�����@m��~�QW�����צ[��+D.�n�C�����s	0 ��1q��P��}�W�0�g�H�ɕw�Z*A�ql��Y�w��7�_mj�cQ��-��}m���|ｑ�C�q����ޓh܎��P���<fC�P��z 2r���"��IUY� �Hz���%fnYW������㯺�H㷧]���9#|a��� 	�`�7"�q�i���:|Il����|�������w���#��pQ�P1bBvR����ݞQ��wz�9�����¹�j���ϫ�9��4� ����}�@Q����٧�bJ�,f?�6��� 6����9�OLs���*�'L�Mt���	��Ak�źV�wa�q�uP�ǛQ���a\�_���ڥY��Az&�I�t����v������'{���H:��	�;t�� �
tФҒ����4z~_A��`�=-����~wHt�Ә���+�ݘR��	V%�j���Y�i`UO���Ae~KĀ����I؛&�.��&0��
=B��0��CN����N�O���n��0�zāx>2QP��xb��䳪�ʿ$뤂{�HD%�$�������.� r2�\�6K��(��2_�/GSz���!վ���6��QM@쁫G�;f��!���y^0`�ǫX@i$��(u'���%n����tP-?\?��Ոu-΁U7)���	�_]\������k7����R�W�K� ��S�)f�(9GUE�P�f���miA��Z/��DKxLa\%��:2�(��o�UX~�(�#)=c�G~&P�E��u-ou�U>Ƀ���i�^�)��Q�z��}<3J��O�_4 �'�2|�����W{7�w�k��������Li�}����~�G�Ԏq��ׯ�ީ�C"*��Y�~桭Wca��}��?�zq5_�p��^������7w���̝`iJߎж[����	��6B$Ěor���uߥ<G�N@��[C�ʍ�`�u�j1=���8�\�d�xG�S>��Ps�E��K� ���=�ӗNGnw���G:<Шտ�q��8!h�}慱��n��ӆ��6�ʲ�[£����i��a����\C<�8,`�ȜK�$�+��;*��5�U}q r<�#{��)mkc��LA��V�{|�d5��M���Y��h�	�
�}��
cĜS��
����h_�X#^Ϩ�( ��rIp�7)Ԑ/*���!��[]�e����"g��9��y�ǂ�x�F/8��-Ggq�$��}�l���O󐔐���c�U��T���m��ʴ|X?��p�Ĺ�^�3�:U�T�Q�<m,�>�(�QT9�ii���DZ{w�u� ��]\ԕ$��B	�����d'��Z0�����h�!܉��,,1 ����zOO���v��Xe阌��:�h3Ž��D�����RvI۵�R��.�������0'���KiP�"��[(�	�[`+�xl��� ��X��K��{�Ǹ��oʃ��T��7��@1%,\<0���^� +��� ��M�%�Ӎ��#���I����وgڋji�쾆����텘*���¡aX�p{q�Z�Zҏ��u�>�+#��ab0�e���Ћ�1��G�>sS��u�,(C+?-դ��ߗX�S<Y*�X⚇��D���c)�X4��6��{@v�)�0�u�W5(t���H�Bw͠U�Z�dJ�L;$	�v�n�B_�����բ��,:P�N .e��1�Z�mB��Դ9^?nuQM�#��M����������E�4S��h*��&hPE�<���~����6�x9��~qU�����`1�=6��q��d2�g-F}�<�,��"�9I�A,����u�>cm�s�P-�@�I��̣�r���h>j..'ٿ�xU���%���~*˃8!.r�YOOh7�.�Ξ�`t�y'K��m$�L��V�FЭ���xS�л'���G���`J�0����T*0>�	tٖN7аE�9X��)︖�O��8k��D�N�����9u����3����>>�+B��[?� ��.�P��8\"����SG9��0 �qi �U�жU�'d�it~r�:-�7�ha��������C 7x�fʚW-�S����hn�c<�z*r���څ2��t�j1�؞����s�^��d�����k��9��rB�}tp����O!�S �F�	*t�_���^�ۇ�E�`��TW:Z`�W��N�vp�,)� Um>���S�(��*|ͽJ&��r{���? Aq�4��c��c���I4��	�H7��6QP����j%3W
�E�Ҏ��$���n��b�lrn���O�T�g>w�h�Z�f�n�$`�"�x/����T��~���W�'��V��UG�I5��æ1*P]�8�������_1l�%o��G>��ζ)bi�ͽuwhR'�قz�z2��SY��O6>ot:��X�=���x��M�������Y0Ҥ� �/�;�+�Ҕ-{-��˧'����)a�P�s���	����$��&Lf�s�͸��7Ʃf��=�Z%/@�������>�I*��j&�W����Z������(|�����=����Mؓ��+�P��i�9��n����Z�þn]�$�y��,�	���Ȅ�3t#�����[BdŇ���8!���C��������>�
x_w�H�Ɓ<����`���������p��D0o�s`����.&�Dd?9]�|R�(�A�0o�¬�{�S1ۗ�م2T�j�6�D!؇V��9$�
��!��o��n6M� ���WRJ̾<��=B�M�2��^��a�o�`��;��$�X~I�(�b����x�>��Y�f��P,a�Κ�b��z�GY%.�U���S<=�/�R��G|)��|�<�dq1�b-��=ҕ��Wϼ���9*0
dI�W��W@*b���y�=�3��R ��Eo�4�y=������&E���iA�6��(TV6��9�3�©�UJzy���?W�o��o��Uxa!fB'�N�~濒 ��M����~S��S���S��̌:v��6��I4V�"��gL��Gc)4`���fF�s	�Ը�'w:�=$q�X�_Q5ۧc���B>W؀��̗�f,=eC��(g=���N���
����ߧL1
 �%_�C?Nk�_�7�QH��!�����J�WS�ؐ��?�+?,i��JM[+�l�-�#���YoW��E*��b6�0���^�G8��D������� �����#� �����Ӥ��s�6/�6M�_:���]�h��H1
�6/%}�
��˗E�6!#�MGB`���@#�G� :ϋ��2&a�P�YK[eј<�����
�����Y����w�d=&]3V��S�҂}jS�*��%>�!�/A�3:�=�f[�)<)[����8W�6O��P���,�7����y�'5d��H�`:��P�,a��51���볬��,s�C���Z'^Fݎ{�FR��b�������X��p4?��ڗ��z[ݛ�ؕ�<�X��IS-�,ω�~qgvE�� 1����s�U��/�F����U��@|�Ke�]1�Z���;.}íq@����M�}��#�?�t��M�OP�	�h@7LܟH���9¥ bx��|;��֍o�9�6;	�\�#Y�r.�1R>y>�N��r�0Ro���D;��G���{v���߉�����.���Tk�f�,KCl< $����D��kgz��^��VN��hY�D/�z�6�)O�/��������A2vjX���p�%��脆� ��W�"N�aY�#����T�b8��	`t�<�7��@�*gWDŝ�}�0�_#A�'����"y���x�)�,'ۨ7��gˎFf������C
��,/{��H��4:��H� ���,�2�6�V{ ;K\�;l��$���C�'�>/��9v��'-�)�QiZa��v좉ʃ_9M^��1�Y�^�Ǣ���U/T$aU�����Lq?:8SGoD.ʋ}.�OLT���0fx�+D�6��<Tá�Z���.�&�[�@Vi�x��Z�-j�~D�%�8�Ƙ�D#p�_���MPi3���e�p	�k׉vX�.ĤlF�v�a���V����U��჊�M��X5 �׎�B.OWy�%)�[ߐO0�/ƶ�Ÿ?��x�����_���@&t�� g����[����>_pQj��Y{c"
t�& "ϖ*�@�3�~�%��y~�43�9��w��8c���m]wŞ�0�t��Ort ��\��!#��>���6Sj�v�w���WG��~��R�Yp^�*��7l����`�Y'q��j�V�a���G{��$.GzЉn<��\��mo?�%͔����p����^C�0[%_J-�f6d��7QU��A����VYZ�R����6E�+f�h��(u�n�����a�H�P����D�8(MJ�$JM�ʪ0�yhtw�w�6�T���y�����;�wK;�ԢW�Pi����б����I�<&�:u 33T����`{�kQ�1�Y�V�k5/�Z&�@�����,L�����np�!b{��1d]�4��o����EvD�)ܷ$��*=�}���0_x�1;Pu�m�g-f�?s.��v�F	���W��KI$��]o�\,��w�Qtb���	U�=�pz����^Bw���٘<�+6!2�
e�ȅl1(6���ˤ�|:�3��mwm����c�����k_*�t��e��k�����J��
+%DYl���X��KfeN��o1�Q�oGwS�q~
����W��[�L`���O��Ss��R^���R5z�ֆ'ū�Z�E�>���d���xYs�i�%
0q˛�����a|0�y������^��h���d̎�9Սx{�U�y�f��?�Vk�b�]��a�E���0�����>Rּ�r���]��[?/0���!�ѳ5a����Os�Կ2з��\��I3�hrP6�s,�m�0+���E��A��	D��k
TWaٙV�0��pk��2����]���������"`�j�h��1.�/z�OT�!��cu�q{[� �.��eQz�`��Lp��[=(�r���tU�����f��\���ߕ�4�����(��������$<�����~�n�9�ca#\�V���ڜ�u��U�y���0��Q
�Q����-���f����G�����k2U��Q3�-��xi��aVN����Oi"���K�� 7�ѽ����5w��(�I)�{�?C�?Q������gN�ˬ��1Bhy��M�pA+W�t����^_������\��b9����gs]O�76'<��;�U��-PA�ޖ���LJԭ�����F�jA���0Ȳ*�,��
1o�jv2B�s���e˶E�>�$������S�s#�S>��9������B�'o_4%9��I�I���eH���t�kx���(4#a�=�YC�X��5��űi���K�hWB[�����K�kuϤ!|ml?��{k.|�s�/�򅟘��f��AV(�L���s[��<I�L�|���θ���!�sed�.�$]ja�Y3:�E7����r1����Ga�%3���~�\eKzZ����-�}ĩS^qC7�rv������%�q����n��5'��v�z�_M���l���3=_C�l���'(M��aW:�iM�]�qLn '�&�\�O�c��y��olt\�/4@�q�q��kC���:AA1���&����9#C4l�N�<v����#����xL�����RBXe$��?S�!��n����B�S���s��m�U��pY�z9�vA�������2����[�G��߇r��]%��Q;{k�m��((��w9�_āV�XN- �> O���lb7���ڌ�Q�@r�9`u���N|�G��b�@�
��T�17���_�|��?R�l����	��W%L�(�)�T�{JJk����.��)�Za�� c���0cã�'�r�X��H�M;�Vk!����n���@sZ-����87RR�M�K,a��1��}�J5��~�v�J�_�֥;82і;|��*MV)�������oiu���#ܱ;��D�X>���?��3��mꘓ�Ǜ�L���0�� 8��I��ox���gqQs�������z��p�*.�ZJO��6�|A �O��&�y���o��34ٵL�w���5"�Yأz��\�/m�@�t.oɛ���:!qc��^��1w�&��rD�T�"�Pӆ#+,���]X�m���֎P��c����$ }e8�]�=�qx��E��; AW�;��N>�����
	��HXA����+r8�.i���ͺF��|(�)���͆@�8�p�!l|�� ��f��]����EGa	�ǆx���7(�-��P�3��.��ރ�H�4-����|*J���v��M� ���G�j6�D`��`���!D�u�]�,TT�����p��?�s�/�T�����+Y_��������]�-2kx�M�͟�~N2B�Hj7�1���:\�> �7쥥����F0S��P�	�㤷��aΦ�|�/>��� v�µ��9w:Jw#;݄z� �K��;N�FrH{���Y��F��3X��(�$�ƗY!U�]�I��,�V��b�����	�C����/y޸>wG�Mp�w���H?���NS�_�`<�sG�U��b0"����z!��	.8�N|�5�Y^�����7Y��8]����
��ܧ�ˣ��o5���ǂ�N ���x�+����ۼ�
y,���Mӂ.?��v�4?�i�;ظn���!T��"����Z�(]L���|�,t�Wh�#�5O�V�	tA�U{i��2#q��ZE�w\�AB���Y��_.��L�f9�A3��(Y;|��0>��O""q�/����}nB��A�[��O�F��_�S�j��|�Q�/[[�A*9ʠ�,RR����a	�T�
��=��w	W�9�>�TĦ�gQ&�ܛ7�w�1�~f(��|W��-'	�M変��r��1��<�pj�\��:�4��}w����.y�R�b`�����$(�].F�ڼ�l��0�`�ޠ��ۻ7	��4{i%�v���Q���D�j�e[-�Ԡb~h�қ�"�L���Wk�e�Ǿ��?���X>�����qi�ŕ�u�L�!K%|ݭ�'D"�����h�?�;)�_R�^�e)�[��Fg�v�{V������3�g�h���������Z���C��Lj�i���=��X��&�e�o�Z7N�X��������u:HA�e{),�T���^ɹ~�oAk�5#V�f�T�^��9�WV��2��Z�p�'_R$�K��"DnV+�?�rn2�E\mhX�MҘW��{�/�
�f=���t>S�<@{W��D%%J�Ek���B덫e���o�N���JR�??�!�B���'l(�9�κ�x3�7Q3Q�d�����*�}�2(1*���V;r���F��\�;|%JU��L�↰��|�C��ks}�����������S+����Љ���h�Q��`_�G�����<�5�Z��z(KT� ��
98��,I���tJ�������/�@�t(N׉��ݹt`T��~>�jpca3UลnZ	�C���m�&B��Nr��2s��Bt�?h��>�oX�[W��3�� ��!�����P4��.A�	T�g�z��-�c��#�i�	�	"�L������,�"C+VBǫ��z����@�st3MmEߘ	�|	�Q�dʑ�c��f���>�����ê$�V0U�G�g7�g�׹hPϐ��dL���y,��D%�>~+!a	�{$��-a�D�V��ui����2'�L�P�MYao��O��G�[��5|ݡ7���c.�PE��H�r�k��J���D������.*�g��o�,��F਌���M��r��u��-+� �yeA��2�2e�a<3?ݮ�̂0��6�Li%�Cl�������;R9(d�biS]���{Q���0�(,c,J��᳨�Sσ���3Qei��V�!ݡ��f�9$Ċe�i9_w��� uR�%>��Y�%�a����!m	xo�'ݤсۡ��ͽT3m3%��t��,���<E#�4��� �Af?0�z'�]��]���Q��8>�h�š���%x*�;R�H-��vP?Q��4nu&��jPET�KE3��I��^-�w-M3��|_dϭeBx�?0v��9�x��dDG<�`r5M�7�ݽT�
҂P�Q�a�S�E��g�e�=�`���{娅��B���[��g-I�	Z�����Ԟ=;�=kßF�'��9�揯/�ӡĮ��#�������WQJhTFbi�¸X�|y3Šp��Nx������B��&Ea�]2\�V�3NΠ6�,ή:�/��� �k���%lZ�Y���o�9�ن��$�2G��4���j$��2(��+��/��X#Q3���2Y���_��b���yE��'��ڞ$V`qL	%��&s0e�H��CU��<�$�d������-Cp7�T���}dA!�F+-��*O�h������_�Wu�O��<���T5}�c��a���g��8��:�� g��}U�G&����Y�6G��^Y�sD�M�M,h�58�)Ti�����c�F�����!�lRQ���y�� ��5��[��"#Ʋ��=�#b�ӟ557
(鯸�tꋖ��� �Qn'q��8�A�4Z�=�9�t�h�%0���K3���P���G��Z������Xɧ0�d��!:ְ�SV�����G>�Rc�M�H%^����ſ@�q �7b�'=���D��QI��HI�)3.�Uxh!p]�<%iH���d���^�*�L5A��΂�ɸS�	>Z��Ԉ,�A��U���wPI�C�DJ%�{gȑ�-���жf��_5}R;<�f���}�b�HY�X�zS��pf���Ή�	��nLp���K�P���0nM�oxA<��:��ܝ�0�$�0���ު�;�}˯�$F��S�H���2)< ���`(Re�(�
�����9���o��6�1�"�}hf����Tkx�<�W��~�w6f-� 01O�n��B��Q�w@�,�����)��9T����^�ɠ��xxEE����E�R�&��Cp�'�2������'_,����m��VÇ׀Ϯ�N�y`L���go!���DRo�nE�ao��6#��V�w��~~�j�j�ZG���f)z*v��O�|��T7��f�aC_b���+m~��C��HI^�.Ӷ���tX����s;T������kC�h��p����
���У��ʃzƻ ��S�"��979�jYY2ߞ ����jLR[�@fa�@;��o|f8ӈ`'�uz���ϯ�W������T�n�Ʌ��kE4=Un��ƺ��p�O�(�;�Jy�� �^&t}h��3B:6��y�Z_��Λe�����= Kp�ͼ� P,��bK~
�yň��jA���tKu�+Wr'�M�6GT�?��*�p�X���ʁ�]�=:�"]Gn��`�^�u��r�Er#~`6�i�w����H��6��-���*��OB��ק56��M�!��y�-M�:T��k!�H�]�=�����V�+��1 ��@wA> �ku�����M���� '�H��U�Ҵ۟^d�5����Z.�v=~K����he���P��͎�
�P>P�������iTCa\��h�d�A��0e�X�6�a�)(���S�t+��Yë� ;�mI�<�T�źi�(f����=M���xz�#8�D��{�Y �٥�*���j�0�R���E��U\�H�����(�@�HM�2���I}��đ��X]�^�C�QU�fH��)VoG�*A�g� �r=����/�F���4�!s���l}��o���l^#\7�JAQ�z�wت�~J��P��/���q'��hѐ�ZB����&�|��7]�Y߸���f����|��؊4��#�א��>��Z���O�>��w��_�nC7h���!�ڲg,��S�+J^�l_s���NT�w�B����T��Y���b�����]8�^*M���q%FSX��q��)[�CЇ�fڟ�D��>�!�P�Y�9���ea�<p\w�g|("|��Ho �#KAj�]`��t�m\2�#�2"@�W��bD�C�`��'q���x�����:>���Z*p����a���m�u ؖX��Ԧ������1���3Ƞ̌	߉����qt��HΉA���~!����B��W[)
�g�s]�g��|XjV;w3.�_���+�r� ��(v�.�)�Ԇ�a���W�v�S�ӣ�lS��QF���O�XSOE����9q����Z��k�S����^@�Wߺ:�_H�٨b�L1j�Q�#��X���b6�4���maDV�y ~��!��|^� ׎� �hѱ<c�X�=���YM�3� $��p��J`4�­��*�:D�aQc��s�!M�}'Sk���i)�員ld�obFuwUX���K��a>�.7�ٳv��*��̮Ǆ�L������-��z(��,&:^���e�rWv�Qv��}�T�cpR���ߵ�d(���-���P�O�����>�=r<n�������CMPt��w1<������=�M�Y���2i�����ꌽț\���/:yF(dZi��BoV�\j�J4�d��K�h���Kf�µ쭒]l^�B�=.{d�~���"�ŗ`��]9��ڂ�@M-���1�u���}��^к(�zR��}��f�8�e�#� �=�_g�;�q�A�+���7Z���I-"9���Q��������CT����~8թ����}��E�E���H2oK[?��xo��Z{!�L�ݏ�k[��}.l����XңA�Z�k��U��JфͣA�Fa_B;�R�o�u@r�e_��i@�i��/YB��)E�p#)f�V?�`��}�����!�L*Y��r�Q��4���Es�»�D��&��8 �6��BK���Jȑ��q9U�i@�wC�.��>�.9����nv���m�\p�gGӻ���ި�������qP�"�c��������I�k��o*�@�Ǆ95 ��/֎j ���9�Q��Xɶ#e#b��^�������Ww�-�5ڬ5($}`�K)s$��5�M���f:;y���	yc���L�/���VB��� �'j���$� 
&[�D��Tt]/jeyU�c�������v���ح��p?y��{��,"T-p����7���Ӊ����Bk
lZ¼$�^L���+x=Z��3�PEU
J�jNY�Xb�D:̅,�e?C0�G�JGfE�-R�G�/I/��SZ~�&�ʈ���ҳ#
��G5�W�R�3=?Y�͗0��Pv�L�#V�i-I"�4�;KWޝ�q
��*�uQ���4%���c�0���}����G1ڤb��'�,��a�;��Ђ��j�TEe�h�Z]V`��Z%T��j���'z���~��&	�X��"h�C��*�o(f�R�X����KU��A��⑋�=�(����6'�g�j�������2ݕȟBA��Ļ�y�wd���a/\�B�:��yP�y�?�P�4O]L���������ܻ��ū�o�.��-ɔ1w�1P����ܐО<��^o���Hb��x�r�h��ֽ�Bi��0�2�A���*�%�Z��Țw���ӵN�K֌�r+���H�VL��W��e�jB6(�gG������4fċn2��&�Q�+��r�DԖ�!,�������
�@-3V���E�9�"�P��С�x�R����X�	b��?i���`�	v��d��u�Y���$�.������3��?sQN̛c�q0>L-��asš�Ǎ��Jl�\Z9�Y~(aE-�I����b�D�4��#m?�x�X�D3N�o�/u��ɼ]ȚJ�'�%�f!qN�-��8,Ж�G��X7����ک7��n����+��\n$Z�26�	)_rE��㞟X���MrS�b�?���!U�"
�vŔ1�B��&�һ'm%%OdgI�^�Z @��I �\ϫOX�C~�D�=~�5�M&��G(L&uc �K�+�_kIfp��gin�p���WD9��Q"-��S=7��@(�
���
���8:��t����]33��-��ot��
^�
�!��_8�X$�t|?/�Ӹôz�� /,{_�%��N���ayƖ��/�N����I8�ʳ�A�@��OoSԏ��E,����u�q*@,�̸�r�a����hU|��S���q�=�|����ߐ�$���%EZ��*���#�<��3tϕ���3�/T�DQ������؄����V��BA��8=i�� G�D�i4&��"Fi��a�0�O�w��ǁF�s?��7��d�����N�̯�]�q�r��HOV�w؇P�e���f�������0��W	nYD��K�5�����G��>tz����L��T�s/�+)�vjO}�,��p��9�b�����K�6J	@vW������x��3�"#�4$
(�g��;P���Q)����{g��ks���{��ؒ�w�;�|�"��y	ɞq��d�#��Vl[�m�N�>�vs{�*���)>p��W3��S}�0��g�r������>��|h���_a�e\Fd_�����,����JU�������r��_��vjH>��x��mڔ�k�� �vYy]��N+׮"����l�WR�6�,�����[bXH��m {�f��!���.9�������n5�T�[^���޳@�(>]S�[��O��@��:=��}c�y�Ӌ���{8ĸ�����8_����E E�4�<Y46ܧ��7���B���*
4�!~����o��K�xĺjz���-=��$�_Rř�H$��@�N*_�y�2ES��љJ*Ц�<�f��궸�(��;��5���oIJ�>F/6�VÚ�9'��x��!�0��1'�*�G$;�@t0]@�4z'u���[c���"N���;6}j�pǔl��w��MG��-�(Qk�و�ڦG��t�5l�pP~����c���Ѣ�	����_!�~P�	
W}�z�_�ѽ����������0%��^҇���BZ��t�T�H����a�1���^� Ȯ��u�1x4)�G�25=*�2߃�;�n�
�Q�]�����G�O���X-<���K�i۠���SDEkL�-epu2�k���bx��P��m�U��۾���`�^�e&=��K�����a܇E���W�Ǿ~��g�q5���;0��S����M;�X�;�c�)�%^�;����7�������-t��<�iڗ�������)��=���ģ�X*7�g]R<���D��O�WU�
c�����le2�,���7q_��I"�����Ld�s\�in��s�u��0Y�����Yn�'�܇Ԭ"c1�텻�V�N�rs���4Q>��3�eW:��e�t�����]NIL$��?��C�X	�l�86S{�9S��%�Z�BX:�"`���*ٛV7�#B@ޞ}S8�K�m�u(��)b���|�"�Y�v���7Z:��(C�hp��2�L��{�͡\�O����t���W��v�Ȁ;?��hW�\�vw&H���H}b�J�3�9:KKf&%�65;6���B)yv�˲S* e�6��7ǣI���7���Pp�yis��Z�X�EAVv��fu��`�œ)'+,˒����E#��'�J�Dݾe�C�:{�W���Z�g�n��wxͱ�U֫o����)#t�PSLw|�&��2	ax�}����h�]:������g㸑NL�O�%?U�\" Y�aB- �H���{n�����mb.����A��%y��#�.��ذk��@�#"�����`a�X6=bDӥ�V陃Ő�G2�b@��9���!K��並�C�.B)�۵��5Tb<L��Q�-���?I���5���A�1yC�L����h��:�ic�
Q���CX?1�t�Qy�����rKԍOr%l��������۴����P�Ʃ@�!ұ��$.B��xp,�gC��B��߂����^��˂o��%�W��ۓ�F�Mw.p.W*�[A�� �.�D���_���[��+��Сޡ0뢝_{�{;NH+-�	��I���,��nZс4k�ܺb��sk�م�3����3�<u��Ș�aH'A�gY��rէW��C��R
�'�:7��M=dj�\T'����
%�w����N���3SKV���D�s*7j ���E�\Y���M�1�^]-�g/C��ԙ�s˸�Į�)���ˬ1&�ӪX7)|½�j�y\����i�Gqo /P㾘P�hNOc��wuT3��i���+�r��aW~�������8s{�R�׬�%���x�q����9�ԣ���{���U|�
�/6���~��s|�\=x�8&�14O��$��R��������?Z�^5�����x���E� �6/�4�g�p�`�o���f��_���!Z�2J�Oo|:v����XR����hI�<L����Η�T0&E�)nǨ�j���s��K��L^$�^/�^����=q����2g��Ā��Џ�vm�a��ْr��k�{�D�)��EySܬ��TU)`M:me��R�pE�t@�b�-�Ƙ��x��'
Ӂn�9Ld�����J: ������ ����`�}6��@���}5V��]t�Dv�A�-�lL%�i��Y=PR���?y�#�p;}�\��������p!�E;�ar܇r^������M��`_|	�zQ;�v�t�9l��6M� ���J�b�OQ�h��VVf�K�;�t�3�����~��>fM{`[^%j�H*4GŻP�k�t�b�_�M-Rr`|y�҈�D�m�{-T�d5x{.��E�%�0]��!^�rc٘���#<15�7N�8��;��i��=Tc��W�	 "�9\�| H��ӵ��7��i;��|���b'��{��U+M '�D9��>Q���f�
��3�D�N(�pͦ��䷧֥ �K�cv�M�L)�W�(G�@�M�h�|����a�0��+���!�:��@��#F�K�U�NÐM��Q�&G�s^���>7�s�q�hM7d�T�>5��>q��:�1I�� p�
BX�e}5�������f��k3.���OS<��3��
��s!uH ���@[���r'|�n̒�������ڗmk\��q'��AXߺ&Ǒ��cI'`1��:+V�W��6֍Ĩ9<�1��i~�1��Kjljd��j�p���")gPo�x4.x �h�1F �(Tq_�tj
�
��jN�ҲF�$���&�O��1�zO���Y���+\�g��B=��d�R��g@E(��9�uܑ9�\b���� �֜�}?����ˊ�i�:2@2�%`����x�5�l?F�� 
?���I-�s�r�3B�Z��v�����f���hlהM����������&�E���y�^��#����-� /������6-k�5�$��q�*�s+���{�}�a;�Bu��: 3��i���0�i�0�\,&�K�'�jMY(��s*r�}˖�@����M-K���9��
���֏��4�g۲�M���n�"�H��^0�ڔ�QG�#�wU�I����Ÿ��q���}�d�vє�*<�Q=
�-� ����s��5bmTִ[D�+�U�oto�.�#�GF&%������F�;A���'el؁lՓ����Tpמ�JՑӋ_�����m����ޖ0�s�f"&����"�m4*5����������O�ۣ�	B�u�.�b�d���-ʍ����t�2����d���O�(�{�ks������Q�T�����)��R��&0���P�;�*�#��x(����b\��߻�t���a�@���O�3��TF#٣�"9o���؂\�k1la�'Y�i	�fߺBܬ"�JQ�hg	1r�f@^�Ls���	��~C������U|��|$q�_��~S�y���clhl�x�|���F�6 ڙ��\Oҍ}��c]���M9���Eϭ���z^�_T� ғ<�~;��L����B:�0Q��&����zvŐP~<����n)�7��#@���%y=���p�,��}���s�۠���>�L��	/��R*���	pnA=�}y�Nt�"��L�R=丮��a�5?R��ns�/D��
�i���=��n3�0�$���b�~��>���V�X ���5������[��*I�
"��l�s� �D��FxNY'�ڎ�E��+���m�9Jc�@B{�1͵�����<��J��J�%�|ew�Q���kk�0Y�S���=��NeRxEM��,����E��,?U~߹+]'�h:���@�&��ҋ�\��_�S�~�#fFQ��Vŷh�?u�ğ��nQ�gFg� ˴Ǧ��Sal�0�crUN҉���o�x��v�}�<�7���%�Z!��종v?���A�y$���,�����ϰ���*������yњ�]*53���\p�y]���b{i��[�ܤI�o|%��x�}���a����8}Q�)QxK��d:�ϸ�@&/ۭƪ+4{��y6!������nǢkLw=:N� 3�|0��!�;��&	R�/N��l�KR�RK��+=���1n>������Pb�R����~�%x�� ��6�!1Ka�+�O¦�8$b��a��i�0"!,=S;����v��7S���u��Jz<�L����'�������7�W��Kw�z*kq�0�����b�Pr�X S�O@wU|ƻel"%�J��G"�¹�!��,��"���>�����@���5�A �v��쇃UE+.�J�v�g ����e�$��.�
Of�Di/+����K"�~|-�Gd�������bT)0^�����u�J}�5Jk���-�S_r���$'��r,VJ
�N�nA�E$�E9���V�s]N��$;�C���S�z;RM��w<�w7
}Uo��l����V�|���-�co����^��S]`F�Z��Lo���'#���G��m_�i(�V�A�juV�i4��f�
���2*@k��"Fj`�_R���Tl,����F�17��T�޸M{K���O�[��?���pq�Af.�4Ȅ��`��y����+�u�#*����i�;4[��T��L@|�m�g|Qk: r��?�g��9ʺ1
fg�}��ַ��_[c��F<�	J��9�?4y���0^'����;ޝ^�z/� (/���,"+�]K,�+,��9B��k����Qق�뫭)c��rn���
S�����l�1����[�����[ܱ�(�OL>�w��zk�N:_D1�N������n����V#a�<I1�a(��eXV��U�"��aK�7����E�0��9:��D���R�]����a��i���,�E��1	�˘��%��d�'?ЊЎ\&��W[9j
65:uX��a��\��j���|���������vA���xL ^�;�E�L��o��_�

�4��4��p[�z��t�nZ�t����7�*;�}�KS9K��l�
2`�FXj��dw=����a�D���}��x��AgF��խ�X/:E�vs!��3�Y��5��؇q�7,���>i#/����	kmU�x�)ף��G���|p�H0f���C�O%|K�,g:��E
�d��l�v���� )V�0]M���P�����o[����<^�^N���Z���ڲ/�o�lx�j�[9�GLge
f��]��␮�Ez/���D�/���Sz���)\�Q�o�I�{c��{�7���pI���҄*��f��t5ǀ�����Y�Ir��o
��C��n��v��H]K{�_�|&}�|���5�l�Bz99�
X�[:-��˶ѵ���뜒�	�EV,���W��;2?��\3�2	"蕮NuҹG�5��%i��j�6�.B����^1v�?ܷ�sϟ���"ʵ��kv�$������MM׷�Q?M�͙�������22��Y�D�4dFR��Q)k��������,bu��a��3�ɩyާ�����u���y�׾iک�3�	��$H/E+��;XJ[|�?�Z[�,G�qj0�]B���$w��h[TD\�i�a�[�S�=���`��z�fq
P���6'-sX�R�I������ ��fA0����0�՚���7������md�q��%�;oO��v�Qq;�� ��tF�H,�h�+��5IoD�GE�"VD����p� <���&iū�m�G����}cM�,��O�ʞ��J�!�V�ZbM�"��]0�H�2L�6�:�Y�F^��<eq��\˲'CD�HR���=	�B_Aه��/>ei���{k�����D���sl�5<蔂'�����-!���D�X���)���y��M�N\d�d�+���E��!	ک� ��?��m7�y��|LV ,O�6�ook�~L	�p���$	�J���3����ís��8�b8Rn_�(��Lg<@��2�m��d��@�{K-�@��K���Q�J?p쥏��}�H���.�l B�z�4o_��s�b�'ui������M�2�r�Ӻv.+ç��H�V�����q>� ��
�<�x�m��Ct�.RN�1p���uqYm�%���M��6%�B/�z��6i-Ƹ{�������&�4�a)��.E��X�0z��(	��z����{��4�fy]�?-���:�w��{v�σ�h�i.ÍмP��%���З�f�R�c8�ۏr����1;Ѫ��G�T`���YOu�$K��� �X_qx-� ^��Cb���VaW���Q�T�)�d���T�����;_ ��m2���X����$��	M	�ȯ�/�$i&�r<�z�� ����r[��	��$�վ_���k�_����t(a�͐}��V����P��se����q�gϠBKNzaOqP�9�6m��H�u0����yIb���z��G�=
�(��D4d���_	<��B]a�Tm�L�d�_�{j��v�DK#��l�6����;����mҊJ �AŅQǇ���2#�!���u���u��t����Ɔ����<iM��.���	�4�,d�/ {����	}�rO1-f�IKh�hg�?jA�����>i�J�[��^-�Uӆ��# �&ں��o�P�\�7�Us->%�Ş��R+3u�:7�ج~�HkC�ӉT�������L����	G�ĊM����Z�wl ����݂��#7/����viz����5��X��t�[
�s�T���	����>x��7jdS�{�r�n40�����D�sq-(i%�?�ʞ��;� �T9����-���qFf���ݾ���=��8��$�ʉ{��S�^Q�̌=�F)C�����n�Pe���m�����W�M�VU��48XVF������Ҳ��0_���4N Qbx*��$���W��e?(\2 tY��EC�թ1�_�a5+�*���Nm)�8�L���CL+�j�%�o��wF�v�D�Ħ�#�.CK��,�Wq����u��7�*��v�������ˊ�w8l�¼Ig�v6�0�[��āEJeQi��t�`Lp�Jn6*WY�;������G#��P���JYzN��J;9����QZ�V�6��i�K����@��+6��j@rb��r80�s^�?}��v�����\�̻�'QăS�Տq��j��uv�j��0L��C���$-���Tx�Z�*P���s��'ui�U���b�����8#*�;0?�eJ��w�� �d���~��o^u:�7�i�����^	׾����h�2�'�@h-���35'���d���ԟ� �-�M���M�L����jT�2~i)
��=~�<�-���{'�A?[֧��5[��O�Sm�(n��K�O �_i�l��'O��KY���E���!�/��YKȃ�����p�A`H"�����NS�l�@|i���u�ϭ!H��~�S��}����i���O��Q�|�-�cH,x��΋xTd�#35��]�9�D�٫e$���NGf�_�80����h�Y~:���)d��F}hq�+a�{Dy=Xk��(kSC�"��V<Nܑ(��/og
��хMw�*�qw�"ǝ��9>���OL#Q�ߝ< +=<s��
>���)�\�,>���LZ��N�ԅ!61'Ã�߮Byn¹�UڀKa��Vq`��
�kJL>"�Gy��	f�w8��q����
7��ђA"Q�bݎ�g�����/dD˹�`X�L�O��Vz��x���E#�&JQ��3���'+K>w�+AO�NGU�������������0ʮU�5$���/aUisI�UkcM8�H�I9{�u"P�!j-E�q׋��Li�vJf�6�q�['<�#-Y��إO�a���ԸN&6�U��B��8axKs��L�/��|1�V�L|��i����H
=�Z�T��]���'�`���)Λ�ުY\JT����P��'���&-{��m�݀8i��x�����b\�1�Qb9Ҡ��<�8�J��^���pq)�f#�G0>��fB�L=.�{��C��R>^��7+M��GG��c���_�c�7�?k�KOL}]��ל�L�<;���Q�\�B�U��a��:*,!#ti� R7"B̑W�2M>���7�u���%�����rأ[�M�Doq�(�jm��E��ԍTćbԻC7M�,� M.��1�2��C�x2�=9��~ �	WHI$�zd���%�Bτ8b�A�XN] Q6j���������2���L����e���M��INi������3�Bb9y�:~K����]C�L����E�J�[�A�ee�eo�ҏD��Ž���p�M3�����G���e�w��*�f7� b�y�!��|�2%G��<[���P����Hu��F�ˬ����M� ӏI��v��|��a��i/��b�JNVF&+�Y���-��-������4��H��jkT�q�M���׫����o�.�e+Ȁ'T��o���H�:4����`[l��z� �Dpl��L�,���6�����N�����3�� 6"���YhS|��������1��ˌ�?��O�O3[�����Y��ɉ<�
��SH�^�ҕ���ndb��V������3�)5p����Ǐ���*9^�?li$��Ȍv���a�U�h�;��t_'s�>��6{@�����o4c�X/ZRh��^3R��{�G�j�m3*˙x���YӬ��n��8:H:�ֻ��Q��-_&-�=o�d8���J���H�D-�"z��^C��(���|�k{�g��� ����a�n���>��dD38`s*�et\%�F��n��G��q_�RH��>z>�'D�~����~0��n�T��=���Opp��g���.�"�W��B�O�b�	�����=< �Wٳ�H̬�y��'AM��+�l��r?Y�#!�Ũ��-���UD�Q�Pq�υ9��[h�#�͒��Q|�q�F�jG<*��K
�8�H�vA�2ģm��Ŭu�]��c�fϴn��e葠���i�bi�yN7FF'@<蔉�5�-�%��Z@J���2���n~�����{��_��:*�.��M�=�+��E���H{9��]*�暅��^ ��X�gYI�	�9��H� (C�i��?����-e�KpOS�Gd���{>�d抜]G��������y0���%�� �ԶC�(��Q��$z2���M5��sa`��F�A��\�5�Xi�T�9&dG�Ul{<���g��^zRܑ��.G���A��*����+�}�U�Ln(3�D�vZ������$����'et�fxҪQ'&�O�>���sFD9��!O�-*�L@��n�4�����h��1�lO9c_��=�,a�#�E�#^}�+���6>�'�p h�k��9��p���	�K���_k��_Ƙ���k��re�,i�O��26�#��Nj� �1��X�Z��T����(\�H����&���(�۫r�.�zx�]I�Eρ�����Fߦ�%�	<��(��N�gu���L�Q��S|Y�t[��[as\���M3>[h&&����9�7v�4�<>��nn�`w��Z��b;>?��q���X�Sn)�k��]l�^_�E�١�8�`r5y�X�^Y��"[�f	�s6NFAVX��=- E ��q�ò�wx[��H�����8j*�V} ��ש	��Io��0�����"+���>��\s��9|��u�_.� �>\��&�;�������t�0p�ak�%�Z몀��7Сq�H±9s���+����Rd�&��-��#��.�BOC�G��Axi�f@W[�� !�;�Z�DҮȦ�s �9�j����3��<�^�C�g�������0��Po�?	��j�����@�킳������m��w�f[�I�~}���־�(ee�L���,u�Rc������(7�{P.�Zx�V�����`�Z0�{�ﳃ�BO���(6�A8? |U�.�u��p^^
��s�5;3�gᄤky~W��/"�1�S6��g��y�k%�@��=�#��@��]�k�sa��
X^qG�h����T�)L��q��	�L�c�e����j�ps@3��Q�쓄#TZB�5� &1��ty���tL��~%���( ^�j����8��X�4�R���Y#ӎTÇo����O�\���^&���*��V����5R��i��9Rp덾u���������~�}����
� ��/�/��]F�J����yɖЇ�&y�x�I!�d��L�K�6�ZJ3�o}��Y.o����iē2�v��P��?&@H���n��ߕI=E���dm���N&�MAM`͉�b�R���P�|��KP�O�Gi^9�;����7�����%((�AbA���5ޝv'4�<Gf)R�^��E?�1Fr|�zr(�+�Al3����Z��!��N=��肄)���I�M�+�W?�	�*P�+"l�m`rm��5X$nOO��2f�Lԝ>�2�N:�);�F��˸�E:�����ڻp"o�N/k�(m��,��@�j�y0g4�Ma�rIB�/@_
�OԈ��V�b�ǒ�?R��^ �'���y�u���@-=s�'�r��CWX`�i�@ �p��KUYg���S�E�m��ߗ���=���7�+BV���K�g�/؛�����Ñ}�Q5�7њ�83��V_���7��1$�w�0�P04�^C�+b9�	�E���</6��c�nFd�.8��(=>k�&�~KN.�eE®z��9B	�D���,?}XIR�d2$#7Mq�S����ӆs��Ҭ�R���KG)x�p�P&�|c���N �Y�(��|��,���`��E�D.0�5��nv�����[!�w�Ē��C���Z�ao�[���rv[�+�/�&w�]7�JH���|��#�?{.S�-���bE� �jN�_��u+ɀ$��o�j�ɮr�R.��S�R�����x�
�?�̏�H*Pb�Ly�����Rӕݷ�b�9��48�$��~]�p��Kg)n�~Ǎ�<w.�A�G����]G���a�J+��;@¼݅u40��ӑ��O�� .܅���V�J��
t�TgF["�%����s���h
�m�ѵ1�6��?��4r�A���^�=��S��i�`4�A�����|�<�����P�(mh]�� }U�g0�_&4�2`;�C	���N��2���4?E<b�$4��  蜡�j���n	[�x�O�Om��:8z ˟Z�v�VR8��p�ˇͰ*����b�@'�X%%Ї�,�OZ��h$�E��n��j[:ǰ�F����΄��7�ȿi��D�7�K�1^�4M�>d&&SM#p�!��v�{��d�If�Vs�GE�a��9��F:�z-5��>o���JpS�b����?*�um�G��Ix�))����<G��{)gL��� �~�]/����<~���ё�;��LJ0��
�[c�|��P
q�ブ>A�L�*C�l�b�\x���s����ypQ�H'¦�e����#djѬ�m���V���EjKxP�]�+`)��c����_�!����bP�ީ��S2x�E��Z�Z�v���P������msa�=��R�j+4F=�s;�N��}���m���:&���Br]��9���7Ou��Cm:�h:�ҷ"�� ���V{^�;c��72��#aİ r2@j!��Mv�G��.<I?'�t�n#�#��8����3��D�5+7�=�������[eeL���ūw9��V�����[��>�ӫƸ�3�����6���z�u���|a��C֊�۾ed�q'\_'�!�8��Ttd�!�>��w��H�O `Ì�K�)�x��z�<���l�x�|�����tw��REOy��|�����?Ԟ7�(�qqZ�D!� �-�md��i\�|RY���6���OjEDI�(��ܺ�t�O���I���PV �3�O<�!'����C1���f�U��,�OB�Yy*����8;BC1�ʃ*<���n���ۘ�Gc>K��C!g_~�rr7���k�d�K���	|�WB`m��@�Gџ�C��B�.�	wu�ʨ`\0+�J��|�a#�u���1����SNu�Mp�qp����AA{TOҶ-��'��`\�҆���jm|m$^4��嚞�J�S�)U�F��ɕ�H-;��*��ۡ)�#���e)�՝+B�Yw=�&SRl�ȃAV,�H�3�3|��_c DL��S�Ũƚ)�h"=9��(�\R�@[1J�S����(�绽;�-�$���Ag�_/��"�CJId�z�չ�p5d�~�o��hXf�n'�M�̟��-б�Si\e8S�Oj�׼V��Y��d��销��~�c\�?d�;U�U��q[^�4K�%�L�}��$�5��I�m�1P�o�j^%O�ƍ�/��(���2n������ZC�fB6�y�\h��t�N$�v�*&��k�mz�;U�}�Z}æ_L:���j?�<_�3`V�L�ŀ� �n��$_��h��a�s����Pk�j� �s-2�|��\�5�����ئ��۹��9a�(v����o4Mu�{��;���V^��y��IS�D�s�H�O�0��AP�X�eB�w6 ��c�� ���f�Ú�Q	~�ԯ����Þ�-��aEn&��������~>���5�1�Ϳ�i�|�ƭ^�;{�6��눀�Q�b����=�j�V|i������[����ֺ8�����q�+j���c�oh���F�.j*��1o"���es!ꢺ=��ʔ���.�Ғ��,�X"�V��)��Y���Kӊ�A�� ���C�h���-�;BV��nq�!�]"�@�b���#��HX�*|r4�����8V�I�����8�6Z�dr�{����0R�C�7Eɱ�Հ4��A��O�Q�r����א��}^5�v�U8$`�I]uʃl4�ߴ�[�w~��4y7lLn/72-�uN��%�<�����16�����v-�-�,�̗�G#̞v ���aY�_�K�Z���J��Cq�j����j�l��VBǔߒ�$�� ��������7����'�0�τ4��!�p����˝K�Lr����2	-�r���٬��\�X�������nF�O��|0"�6�@J����S�w� �7\ zr�}���x�E��&qe��S���T�p3g�k��9�
$���~��ޭ�j�.�����t���AKr2l�%�d���^m��J�;Y7_%?��L�u%`׷�6 =[�	1�ƊȞ crƮQ�%�g]�x�*�9Kޢ��M���)I����Ie�L��LH�cjp�t�����M��|B���$��ˏ����P�.
�Q�qЗz���f�~Beos^ۛH�)��YF<�iI!.�<���No9z�#�i�N~.��c�,�夕����=�v�E�xװ��yd_-vw�kVτ�9��<���E����<�}�3��Z�5�g��P~�-��_�B����P�>�����sϢEX��2}�g��ׄ��I���L�۶�B��{0E>��W��Y��p� �x)Z��JGƸ�S����o'��u�|h����t��-�'�MaPؒh a�7�J�����-��F��".�:X#���	�*x�>�TB!fx{r�h`�R�!B�ds"��]0"4����L�O���xx}��Z��,���0���G��q�Y7#��)�٣Tl��D����Mvj39�.��5�8l3�g�C�Vxھ�\e�3D.�E��:G����ꘆ�ho��A[�c�a�i��W�
����d��	r�A�-2�`� �.���6�b��`L���u}�'ʃӮ���H����3k�-��r��k'�-���o�,^!�z�b���k����>N;z�슚O �#�Kd0I��ʰ*�I��1�����)�>-��c���4T�L�1���^�;����B�XWK�u,-�F����I�RsҔC׍,���gU-��ڝ�b��ZO���t�#˿� �F�����j�[X�=5�(Э��_M�D��x˰;�ژ�3ͭ�Yq��3 ���VOs5��J����T��	:����[Z��J��o��#�x��L ����0/�$�H�D�T*BZ���S���z�א=��#l ��e8Po���������9����;�������H��R.9{�ӣ3W�|0�c'M�`���K�q�L΁o�jiϠ�W���`E� S�6�h� �z�Z�����?z�8����4>K,��)��i�o� ���?�K�e�� ��.%�m�W4�zv��ݷXB��Ǻ� {�eČ����n���_��5-��-	��N�|*zo�C�����:t2w'υ�K��й�t�j��x[�*Ɠ���x�����������Ң�W�WБAv���,:�ҹ}���x�����˂%�O�Tm�Ѯ�O4��ty���j(��Y�0��q�2z�V�:ʶ-S�f�ȟ�_BC�����OM{�P(e�l:#���5���y����k�D�xE��H����bX������PP�w�.iV�k��D�d�^nҰ-ˡ`�^c�_���`��-���(o<����F�N�$2g1$[���z�G���6a�AJ^������"c�ң�b��-[�Rko�F#�*�/�!OP��xO��:f|^rm#b����\ l9�z�	�S�ߢ��pb\3 ���:'~XL��V3k�;Э��z)�H���B�Uʩ�Hm*i9z�]��pIȷ+&�Ǯ/�
ע)ÚV-}J&�չ,ߖPn`�"菙��2�m�򈾗Z�{�����_dY�YAK����������3���Ü�?(���e� d�0���7��3@[�F��V��	�&i������[
��v�q%�S��c��&>��7�z��6h��p�:�]U�Ą[�Lƛ2��D8b�J��;�d7GSb�Y���j��z�}�(<�3ϰ�ŕ���f2�lv��V�^�p��~�\�~��&��8�{�"L�"������k��!���w��D�<��t�ы	�o�գ��-���?�,��7��1���'{e"@��
��O�~�85\��J�B���Z^S�� �R��˰���+O���m� ��7(40�C ͉��F��p����L@�L=.X	�Q{r��1̳�W�M?�m[�Y��״IzwN�$D�ђ�JF�5����[4�\�n���ŵ|Iq��ֆ���~���>ϐ�gS�x��f����T��r�V�J���Vw��jI9*=A���ko4w�U+����bP�J����+e%J�W��(�=�S���';�5m�N��|��7?F�3��T�ohq�GFFvς��1Rz���+;W?�?����ԛ�i�<?�5�i)-�mTk"�
������7Y^F���'���s����A�悵��R]�C�]�:��NfOc�J �"t9��:Dǒ�����J)nUy��_D��=�o���������߮1*0�FX:˯�c'��[`y«�F3�]gg��A���	���X3	z�)�d�G$�[3:eD0��N�#B�#=#QY�,��ɥEd���k?�����r=&@M3�d4D�ǎ�(�������Í� ྫྷ���k$`�%�&'���)qa��Ar����6x���=�-v��@hз<���,@xHIl�����2�-�yҐ�Z��5-����a¤�l+t�t�0¼��'��0<A�ev*w��X�hnp;�'��s�����"Ck��������0u�sû����k�m�ǔ^Z���� ��S
��]SȂ��YW�i7�^��<�x�jx�C��8Z9��ߜ���K�m5��J�gCR@ x�4�4��R�C�:w��W6�:��Nh��{��q�Ll<?�CV��I�S�1�.��[� VZF�^#�����IRsg	T������/��K�=&���0b��8���
b,����֢ϡv�!fsR�*e]m���0�KyUi�LD�L����~b#h4�L�2�0��JJ�椒Ϥ�4�u�[v���O���Bb����ǒ��ܭ��=��>���A�䬩�^���ivXͧ�[2	t~���]H��ۍl*��~ϋ1^�{g%���H
�(�8 Vr���V�c�d[�!
"�P�ȩ[.U�)�>#rԞ�%6�QEE�[ Xd�����m�	|^�moS��[T�X.���b,	���V�!ཨP����fK�y����}9Ğ����Έ"��b���AB�\�v�G#�a�J�U�Ej��%�Z�$�,�$���1����V������T���ұ^�lK*d��!��J�"�^��X����_�.��������zTz��fbd�06�dރ��|���k����OQ�F~�l��<� 4�~�mPz�Q$�*�5XuE�sH`�5�3R��ݽ̮dq�B@m?Q��y�D�KC�hG�fw�'�"����#L�>GWy����f�|��
�����0�6�%L�S _����.Q���ki׶�<�)LVde�����_7��'��`M6����;�Hz�kac�V�x��lT��*�::a�S|�kd�>�ި?��+���5� ?ik*�ꇭ�qi�D��i���I�	��kO�8bw�߅����Oě����5���h�:U��5��^k6�s�C�1j���;�_����/��fjQ!hd__�W�I����{9�R����I6ěk�L��h��buR�)�%f&��5�;A83,�u�T�¼��uHu�C����4��"�8�2EVx�}w��U[E�?YB����u�z�:4�c�	䁝3~��XN���d��:�a���V�T��h�耨x�	u��� |\ǰ=Y�fr�`0����>��L��n�OZ��VV���4��k�䅣��5_��+
�V�Xn��C����L�X�$��̶c���N�ú�51��u�������
'�%���a��)#LA�|_�Di�}��X�������#�)��k<ɿF3�����P I�Oyw�f��e{ä�8����e]�A��a꠰C�p�SqPDn3n�]�
�zuR8Kl���4iY���}�'J�i�޲�y&����1��I�x�kCJ�	�x���� ���n��03�/�qY<���%��u��p�S��R2u�z]^h,��%������<*I���=a�y �^�m-�x4�J[�DAU��8X(Ҧ�n��0�sI�cC6?�	 O���:��R<�O�A�.j��@�ŷӺ%�.�@�S�(����x�y27��v
�Rsݝ�i�*|���@���_ЫE���8���LV���K�VSn��~	3 "����KJ�(�r1�mNA,ȷS��@l^3ߐ��j;?�[�˚����+�t���'�(��\�l4S��}@�f�/��oG�k	�IT�}ř���'ѯ븆G�-���g!��e���i3�Ky��\�ؓ���l���<�D��!9��`��	uG��*�i}��Ԇs��
kk��S�@1��c��ROl=�Qˆr�6��z�<��W�m�
��� �|���$EXc������|
F-��{�����a�%���I���+� �{ ;C�5G�r�a�XI�zY��W�����s[d��R�^�q` :,�:���qX�����VRض/k/�ϯ� �,N�[�Q�A���b���H�u,��v�[H�8��;0I�}�e$ز��Uܤe4mj�Ψ�z#�4 %[5�~��~#�B�%���v?���Nڡ\[��]4*g�1 u�a�B��$��,3J��������ǜ\�j��0`�K'?�	��Ii&d����Ȋ�S}�ޢ,�O̸pp���ܤ��Ίd\����2#8�(�fÍVe ��1�x�s�󃋜\t����-
;By�q)d�G�"ҫ_��i�?����uz�5�%c2�z���Lսՙ�L��b��u�6�Q���^P�H��S����D��������s�|Ag�%~�T�f��)�� �X�}zʄ�)�r�I�|��^<�W)̫���ţ���J{/�yO�
9��sk��RCy����&��>B���k=I+wQV����%���.���#���O��;��P�F�Џ��p��sOe�=_�\�[����
p�p^�F��>d	5����d�%!ԇk�kyN����A�|���W����x�^�Hc�-�Ha%۳2?a��~���.�;�9�ȩ�d���A����ٛ�t?���x���v��Z��TZ���(7 �t�O�,P�I�qk���H�WR�$��W �B3)��>-=l���p�I�����TD_Z}|)�
�~���ps��3�C{���<;�n�V�Փ�ƃz��Ԍ��M�� �;�4ޏ~��y�=��|�C2��if�-D�!Iq�
jF����U}'��_�E&��f�(�m	��.�F�r�p��^�y��Z�-�#�>Ze^J�J� $�9�6�)Pᙧ	��ߓl���6Ph��$D�c��ĸ�t:����
.w�.��,�B������>g$[���¹�ua4zl/_��!��k ��V�-�Y[�w"wF�N�����֖)ʣ�̈w;"��q�.R�n��	��D�6�@�/D�>ش��6�R�y�J6�@�ʼ�^r;b�L��C������&ksqL���B�N��%��y�un�~?/^a8��M��1(¼�q���jH|����a<SO�}�p���pd`��܊�O ��ٻ������ߐ2Fw�����{4ע$-ϗ�("%�6���r�����&y(1�R'�;L9z���s��_)Ϫ��(h$ڬ��m�4�@�����\�g�	���/������o��j�GC%��ŗ�
e��|��(�)`Aղw��^��F�����n]�����.�N���ۛc�O���Rw�m��LS�o8Xxzd�7 d�l$xs|ې���P��jb�~"�Ю;ō�ƤK$DA�=�,!)⤖[��-W�bOژ�!K�l��wI����<�"i\Ph���@���Ǝ����"pE���c��$D�⛙%T�S�]��*��z��-�m�����`��Q4�EЭ���ܢ4/����;�O����a�Q���H�/��!���K"�������Ekq TB�}���W�(ێǍz���1�h����c�1��!ׁ�o9ܷ��zWSt¤�yGO��w=.M/XT(?p�D����}?��Z *c�*�Or��2�[�!l&�W��V����
��k�g&}�4�Y�Q�g��}��Uk|��g6�?.<-�E�%C�H���� ��Y^Ҕ�RuF,Z��;��VJ�0?Y�H�r�)'�2�8��m��\����_�
=2~�v��As�d[{���c��0il�|k/.����'�ܝ�c�UeFv��0��� ��!!h^[���6�.�l��sh�#_��'(N'r�i+,��֨�R6�lP:����2�e~���Q�r	va��sn����;/Z^s�@w)�鮔��������ܪ�Y��C�ޤv���;�脏H�n�������G�n�/e��_f4	��~{�lx@�(����g���Oy3f�H���U��(� ��_ٗ�ᓭ��%�{P�ġ�r����Ũ�[�&ɮK�I��%:[pF>?<�p��I�:`��W���EU��!7��[c	�CUz���8��{�h�b�}CY��� �S6a �}T�

w�C����l���ψ�4�,�<��W7#�c����|�(�(�Ɍ�q9�	H��L� jrTb�@1H��c4+|wѺ�G$c>�}�:t&{�/�����q�:.1�ц�Q��B�Tv�@&��ºF��	�
�-tJN�+��8��n��W�1�y�7�XD$%f�^��� ������q&�*�����Pcj�x�)
T�c1\/�4b(�:�x�kR����V��Y�-��0� i�A-�y��0:�eK��3�9�/�W�\U'��լ�p"ҕ)��O(��P�M���[�g�h�~�T,*_�(�l��ڼ���ۊ}�jz�x���8�x��>�ऎb ��I@x�M��(|+�-�/���߇^��`�$xd(+�6
۵�h�[+��I�B���1���4x�@�@�| ����Z��2��A��'3�'�Fs*���U
�{��x��H�ZʗzC��h��P6�,B$8���*��+9���ɷ֏��6�X?�\�d/0�L�e�E��P�g�0rw��g�1�!T ����¯`\�Z�#�6W��|�P�U{���(G�����s��XK����	���e��@�y%;!��":�F�����i-��_۵��0 E1���:`y{�(I�� �\L$Iv��hA����<�('P��n*�Xȋ����i�bcj$RA5�� ��~�Dr|s�T������xo4
�_�*2g���aMn��y�H����v��uT����y�����f�W�����z|0��i(/Hc~�ӬŌo��FH��94}���T-�47x��E��J2p��Qt��e��Q��AӉ��dJO����z]��ֹ�D`�u}@�_� ���+����jȡ}�H���wRXV�d�w&1D��/8~_�(Es�+�W��	�q�	vD��,���L�D�2�&_��(9�s�9О�3C��mF�o��q�\@�$�B�7ǀbr��'������h��)�GlN�0n5@����	�s�ΎzǴ�r��G�|�c_���Om�L�c�`�.�8��!ʻ��!�\2��
�!$��ٷ����!T8�ٹ�3���S!Kt<�0n)��[Sm�K)���+�9�m��%�U��U[���0%z�/e��rh3��NrN�f-��������7�,0D�c��L�������J�����;�P�M�����~��IIa���\ګ�.bSA3���	��D'ݧ���UJ�Ntؑ�:]a�;�<�8`N;�i;!r��*�l'һ�+�0�=��|����a\�N�ި�/�y�	B��"�Y)e��������He~�U?�]]AQHS�h!ϗL�$4����r�{�ۇ����/P���}|~\O"�a@���Ĳ��Ї"��9y�I�.'���`�>`��e���yc���
؋%�ɨ��FB4�w���:l9��p����s�@�_։W� �rt�0��sy'��$�L�;2E��d�%雬���Ȯa��@fB�2�c ��a%�ɠ<z՛���&��׶N���#?Ǘ���-�Xy�d}.�
����ǐ�j:�=>�ge�4;�<���`jթo�q�,Z����ݟ1�R�9����rn�!���-.�^�K��l4#��,!!�O�K�s�C�k�����?Ix9¤���nu��*Jl#�B}���ȋ b�c^K7���d�����ĦhF]�oB�)L�<f���O�\|�9B�|'�г�ʘE��}���d.SKΓ�CO��m&�#����+�#|���Do:�BO\����g�?�8��o�I�a" �dӵ'-�*��%�o�e�m��\�%�-�T<�N�����	?���h]�nnM�(&����sf���:��͈�X�H�Ζ֨�@�  I�ɑ�-�&�6������<G��%�{�|b�W�Щ:��&��Im%��f��^>���v����L#ܚW�:���p�~%Y_�����*�'���BFvַℜ)�6k8��+�iL2�Ѻ�pD�	�P~J\��Eޛ����k�2�r��kc�]ǩkf��gl����,x�\AȘ!�t����E�R�R'�ˁ�ݻ�֓a���Rn4fs�F_Ɛ/�ټ��X�;C��ƌ ��]���s4*N�|�RF�@DQŤ�t$���נ(�T*���^�8�|f��a��d:q��R��Y�In�2��ޭ!�촜�T�я��l��~�e�J�)�A���.�I2E銦�+�t�2�y?�t��w�6���4�.�UR��X����ߎ��ة�Ѱ���6gX�6�[�l�}f0X.}X0,��e��X�i�nˀ"�]��s����I�ʗR�{$^�_C�<� �M�BMl��C����u�c�V�΄�0ܧ�{����aW�-:��MOT�v0�y�sP^"�Wt��N�c�!$���8���ϫ�:�(��
i�,H5x��
�I����U9�AM|cn١��g��8��~�H)�crk�c 3/�v��Wyo�&��\��_L��v5�����p�1���wx�5$9No�rZ�%����Ü�%�{}y����ɿ��&�m��x�ˁk��2r��H@�C?D�t��R�a8�G^�^�.#�j��>��4�6x��/[��k��個���'[�46�j،4���_a�z=hYͥ��1�� B�I������T������g �����Rʂ�}њ5K�u@�fMhAs���<y_�S�"]�0R��d���\���i�CZ����$��z⸮���g�Qj�v �ף�D-�be�r��^���;��$([�F�oQ�G����_˹ő�*B�����x�����JW� +�*��W{"�gC���N��
q�i���,��,�h.@�K���,it��*��r.�$7�Z��FEzQ��S�Arz�q5�)_�$6��J���^�g������Ϧ�H�Z!x�bǎn_)�d�����W�А%8}(6�!��lQ>JE�#�?Y~�߯��1@W _�r�lxc.�?dZ>P+��5b���t��얠���p�ng��'�IN�Q̰�CH�aftd�E�:_4V=��kD��.���N;�
J�"��Hf��\���۩4�3�Y�\𹘥z�8��>�`�srDB�<QM���J���}�#�y�1�o��iv�L�%�>n���H?N�@w"�U���V�ݻ�Z֢� y62���U���\.߬P��{�l`oǉ�P1��Y�du� �t�V�10�I���:��d��&�_t�SV�g��B�m�@�7����H��#U��e�_I���g+�e���d� ��ҕ�����D0*HZ%�I��{i���Z.ʕ��q�W�<�F�&���_lɜ}T#FȬ������Ԕ:I���Af0�
*��J;����e0���M��!Zs�B�V �[��[�ށ�/�(y �:i��d���ҩ���ZaF:�ĸ�7zqdF��0���$�7]GjS�@ъ/�))�]��m�[��Ɤ���n��`3�q���j�D��d�\ۉ�8��<8�C�8�����Ċ��M�͹23��X��������D ������
8%|��%�a~
>M�瑈��q�1h�XrN J��nH�����C��OUU�#tZ�76�Dt�v�߮�U8��9b�������ӎ���;9D��sɴ�9�=u 	��*�hx~v���;+��Nm8��(��g��/����2S��CX1������v5���&����<NJ74������v2Hh)���E0j-|@��ʈ)O��g[D�m.�}��J��E���k@����8�#���V���)3��C2p�)ۺ��tK���M�.iG����ח��_�~��z�Kݪ�fm*ا��R �c@���Ԟ�����w�۞�A#�k�:0%���GkG��9G��82?���l"��N?z?f7'c"��.��4^&J[� C��3υz,VU�с�=�R40��o���)�����v�֖H.U�׵����f�D����i[���������G��-���l��K�]�O5�h<�
T:#"Flm�1W/Ӵ��fb��(�����{���V����R�z�f�;�SF�� ��n�H���%�	ۆC�-���\2�27���/��|�
��R��M�P��<o�����:��E���`;6r�+Ť�V��1=��H�����D^���4�J+�4EB'�z5m��f,�	�pMD�û��4E.��^5ձP�"��/�v@�wa��g,H�3�_�'�"��Íd�����W�~!Vh��P""�#��t�<tzC8����UEp���@�O��ؖ�m1�p`��W��,�I��+r'�[C�7H����?+��>�N��T=����S�x���N:��d��I��� ��l�n L�/�]�� Q�<Z��4Rj��C�Ŝ]�G����	-8���<�F�r V_�29pa�N�CuS�}߇��z�Za<��-�c������ݢ6B\�"�\�8NOnun]3����)[؝n�|i���Ȥ�X�;����J�:�A�>x;�-!;������q� ���G�j�Խn��K�.�

X7���80��]wv6�!�;�������P�|g�j䏰_�j/+�f^�+�e��J:JWJ�� l4)��)��&>�GL˳��w����})�)�B�H�*5��?����t�&M�yPs+ia/#G���0T�$kB�e�Z7%��<˄�h����(�����Lw��=���w���	6[d�+c����g�
��¾�����Y�1�1��M	������c�'<����fQc���y���Z� LMOdP�9��2���4B\�Rt^���
�8D��/I�IO~���Gb�Vy�ep�J���N����v���n�w�xqj���}�e��ˌ��0��$K���K	�V5��l[��S�����G��n����Z,7���>-t{EH��86C�;}M
4�(Q�������X�5�v��QQ~b_8\�N������eS��=��̡d�Y�ۭ޵r��<�}�����'�h�^�!��\�p�0x��^�)MR��z�7J�$��D�B��_��[S�n)�ʑ�����*���Y2	/�Dk����IQn9%
Ķ���|��S���pb����&w��ōɊ8��PJ����y�x?F�kB��o���,E�'�6VoՖ1�<�%����"���7�|�yٓ�NM�C���-,14�v c�{|wo�4�bFg���1���f}��!`*�*q +!�RPg"���U1�/<%�{0���9�����x�#��p�1��a��C�}��k>��W>�����r2�>�`!��t!6"�Mml��g�4'\�X!7��<��C��L�~�j_D�W��ԕ[b���6��KX���-b;����37�(e5����x�Q��okxi�Ώ�̺L]�YA�&�� ^�!x��;l��cb�@��lu
�^V��۵w��j���Y�1\W������ ����R8Z���;�p�w��ҧ���Nn���b��ŋ,�c�ݦ���c��*��V�t�f]u�e��4a���,$��ʝ�uvX�: ����Om�'��CV�)��m"`�����#.��U\W�d���^*��2�+�^h�\(2߬��V�sX`1����t�C�^��)Y���dF'�Se=U�2>����<�[.��v'W�'��n��Eo�OW�Q5F+���J5���;���%�8�1q� ��Pa3��D��Cy���;�������{��t���㥓�G�|��S�z��?mAa��,�&�Tu4�W�M`RuYQ�l��Nd�w�V��F��F�W��:����! �$0��"��u���~��o��^^�9������N��r���Q_h�����õ+ul<�?,--�ݳ�f~�2�N�.�,�r�5����9�� TWF�ĭ���@��}�����uk��#Ց��<�K��i����Xi>*1Z�^�<���Ps���H덱Ì��A"��J6�A �?�1;�࿔��!�i���!ot���ZG���xkm�����,�\�x%����BF�i:﻿�	o���ˎ��3�����!�e�H��ѧ��gKi����R�S�;c�^X����T��zHY�5tۦ���F�d�������֔ �����!��?"��]2��_�{���N��w�-	6\,��Z��:�B��Bp减e���2��(Pڼ�x<ws]j�t���
g��JpELn@�/�d�3� w*�F�3Dz���r�
��X�+PV���F8�+�th�͂x;�vR��a /��k[��'B1��j��9 �p�B���s����/"%�aO6��MɃ�r�q�6N�*A�}�~p�Gk��;�59kM�h�kTIp���&w��
^=0eE�B�b��P�X�{Ai߾��}DIrc�B�WN��(l>��ٓ[(��*�(;�u�Ұ��}�֗O�����+��w�ؑ�+O��m�yW�_t�n���:J/C$~��4\�o#?��,��J��"��۰em�2��^�F�����,��cO*7jMv]G����:>���4u�"#Y��R��{̋��O���|��|С��r����.�=Iᢊ/�����T�@����Ŋ�H)�mXC����ƾd-�_�ƹ�<#q�H��jx?*%�%�p#�
m�6]��+���"��n��ڞ<E�Q�m�QŚ��,^܉�������./O���ooVq���
fl����0�Z���]_��0����B�%໣	&^��1���@� ��~^٨w��9RF?m��h�=m���iZ�$�S!��	GF����K�4�5~a�����g�WԻ
�6���X+�t��y%+Kb��m?Ȥ�v��7���8��/mڐgl����z���^SA>��f��e�����@Ԏ��k����������`}�F�_�����!�����!��G��9)O\L����s���+P��Ki]�cW;�D�L�T)s��9r}"325�V���#0쓖��v*��Ba��&Hp}��'˄@+h#�y�FeY~4�g4�\{�5�}���g�OM�!D�h���;�w6Y��E��lj^�/��~F�d}r�[�.*
;�b�7��Tf�	 ��}b�����{!]'��Y�s����bі<����TsөC5�ʏ���1�&�����"��4�y� "��=�?�K�ڵƕ���t��L���W��D��"6���V��d����R��VF�*n�j�ɞ���f`����tNR��.�v{v�F�IVI���4�"oM�r�:�T�=oI�n��i�b�	['=T� O�]�Z;y�smN^�F�p��B4Di��a*�É���&5sT�;D�����0#�|�����9�������O��9���F�s�(S�O����ر������F�Yˎ6�F @)B<���Ӥ5�1�G�+�.X�;Q�x��Z�`"�^8��*f��"d���p��
-�KR+�l�iTr�E�>>���
	��<��y�OF	x�Ex���k��.��7��7}�1V���'#�"��_a<��-ݦȋ���t?-������D�P/�*7d=�݄8��(�.R��ZX��p�9���+}�ud��������<	A����C�<�d!_;Q�u�,a���3��gURR�5)��ύ��
�����MCF���?�Ӑ��C\���6�;U5^X3W�T�-�N�N@���1{΅��p��(�o���K�I��jht���������E�/Pނ��Ѓ9 C��3X�GO���;�����r�2��IK�)oMȗE�8A��0[���4�y(aX�ͼL�[�d���tu���1��'E��<8�J6����).�Ti;@�K�IQï]�"�	�/t�B�G�T5��?��3_ZR�wU���`��Bl��A���棡��)yA�aC$c�6���C�F��ނ05ׯ�^��'����/,���n�3�P������t 7 ���A�I��r�jŃE(\Y�1���9$&]��[����i ˈ��QUʬL�k��	M5Y�TcA��#,�4��+Jq\��D���!bᶎ��a�J5���4oq��|#��!l`*Lk>=�0��n���̌LR4o���s�/����:�}�z�Ɣ�}�����M�c﷠v%���*�
zq��t�tU���W�B�J�x�F��g�����X�.Cm�Q��	|��<�;����{!�gk&�}���&<����'�6F^,�4f�m���㻔Q�FvF�$�i��v���G�jt�j"�=�~���M-S>9��^T
�����vJ�
���I[r	�<d �b�"�+18��p��'Bq��@�J}�+�H���x��ږ��=Et�M��� �?Q,���w�W���89��9�.xB!ngŃ�w�YI0d��5ò�~��H��o���d� ?�rRPq�zL��!��n����6cQ�����⫿'�&U
�ʮy����\~`����a֚JfsͿ�y�;�;�T�7�ML��l�U<�v\:�EQ�'e)�w����7��i�����؃��l����<�B�٦ݿ�/�X�f��U�C&frH�0�na�d��Vf
xb��sH����Œd$���'��)���;|x�q�Li�PC��x�G̒�$v_�'�V��0�^!���1���Z�ݶʛj'�����#}j���g/C��"��i�����w?n�X�L܏{�"P+C�&_tX�w���'�aLif�@�%�Zێ&j"���=g[�Ac�e]�&�БD��[��8֎�j;i��B����e��W�(P8(B,�5=���>���5���A"���7`��-#fdg��G7��rE�I|�3p��ښC7J�㍝.����ٯ��_L�1Ӹ���ґ'P?W�Ȑ�����d�B���o�������ѭ�+��\N���|�Z)ׇ��מM$v}Ԃ{��:]
�	�|�S��6�nj�]/v����ؿy��#���|C�/��U��3��|�NĽ���9r�X���,�`J��
>1v�SQ����=H@���I��oyv[7�X �)�؍��r�J�~����^���e(�BϨt��c�S��w~!��0Zߍ^"�s�c, ���Ǝh
��j�E��G���m�ҩ��l�mÏ��%�$�v��*&�O2��w��!
���~0�Ĝ�,��,����S��#�N��$L=�1�F�g�gh)=!�����-��U�Hx��'#\d]fo��q ^2ڋRePG"��q�YP����?z��<���՛�M�%���
����ݩ�q*��y%���և7�?�B�z"�"�w�s\�Ъ�T;���C)>�*��G�Y��k���W���Tr+�w@|�lۍl�w�A���5��<�xۡk(9N<�A6Р���Uh6�\6䰴��c��{~R�֝"b#R�3�׺Whz��w0I7x�!��#0��S{5P�k�4����u�h`��1(�o��_�zC�zY�$Uls��F����B5*�����5<d��;�)���F��[d�� �d�LHD����)P��ʋu�\u9K�'o���Z�t-Q][�[a�85��A<��F�I��`���zP46�?���]@�ԅ����EJo�q�|ю�G�Ds�Lb�XO͖!�j�@�$�Oյ�R&�y����bֳI��P,��A8�y;v�l���N}֍Y��е�ݛ�]?IE��(]�.�u{�Ȋ�H�p�T�Β���Qڢ{��<�!}�BD%�H	ҟ�n�-��Ek�}db�9C�V�1�.}���j�?#WK�6q��
_sL�/��hF�(A �N�H.�3��I��p�r]�2�TF�C�B9gޤ �Tpn�H8گV��+!F�?szۙ�:V��r�ٯ0��kP!ѧ�ҷ�钫&�G����Hbp8']Q�Qv�6o�U��iA�|ć�k��X[�r�Zf��$�"i_�`o@�[�`5�IѼ�G�6c<ќ����������]��vW*�^ h�Z)r!�-�'>��W��D	�^s��B6;ٚ	�R��W^���B�=�g��mc8��ĔR�?8��h��G����ơ<�Qװ�}�5C]����Mӛ�o���k�ك(�p����j���ou��>yb��MK�5�}�j� ��#�I����m�
"��+lˁS��j�����>����
:�"J:�u��0��.㹇�D �l�������SD��^1R���l8�|���{��A��jeAy��ĝ,�,M<�)�-�����b:�^�
6*��jkB$��~��6	�5���k�ֳ�B=i�uiO�tN��*�%���ױ�@j�:e��"��k3w���b��k�lP�������d�)�y�h�\��Z���{�O��#�=V�(ɹǘR����lڲ�4�^��Z���"]�`z�������R6�%� E��g��s�_Kj7D~J�Y����z�e(2�����К&�͈��P;ZPa��H	�a0�]�1�8�jΔ��n}Zn3�j-����eP	�_&hx��G��M���GyP Haٜ	�O����S	�;����> ���P����^.��z�`�]�R� ��Ԝ��x#:��m  e�[�����*BѠ}
{TD���+�����Q��B��xR������D��1���)���.���V4HH��Z��pD�߈62���R-��t�ǌ�����~����g�����f�SD�ҙ��Y*�r�X�j��@ �d��Ε�J�9�t��|K��)՘_<Ǥ�䥚!���	�ez�J\^�֑�<iwؓ��Kj��6��l����]�q�fy���g�M!8�o�K)y<+�����\B�+�>���Ad�;����9���"I�<��L~(l���_��B�b�5����Ԟw �p�aČ�yi�^�-�#A+��������b��&�u)��!�=0����s��<_��a	Ht]��T����_�Dʊ�}((}Ĩ ���pDO<��~��T~:�t��4�f��?��|'�����t�y��[�~�\������x��^����(��S����{�`�!^p|��B~W��C�VC��v��Q��W�A;�P@׵���	�U����?��@C{�O�.��n�O� '.!o����ʞ�l�^��`����G�!~P��6n�7��u8�=y�����e�Ҧf`�P��1�B��|�ڲ��Wa�oV/�iܴ�H�h>������ʟ񕎒k:5���e��g(�D+,*�� ��F�1��oce�W{�� ��hA�'2)�����SPT�z�q��jJA�/�� ��q?�����E��N�Ш�"k�j���	D�6zDVX�GN	Ŋz���O ~f�!y~{'{`�'U���*�B-�B�%�J���p�˽#�N��h�I���Ca+��f5_#�� 5�5E�݊����O��t%G�;���U�S�v�z9�������������/%$~��)��PU�m����*�u[���:��7����=���|9�ܛ̬�5|V;�3뎵`�*��VYH�d<v7�#J�Rǡ�i�Ct��+f]�I2�Gx�X
�*�����ǖK��**����f��co��
���Mi����I�q��;̊z*�h�TdXі��ұ?��U��x��W埣���MAm�V��M�����W�L(k�E��|��_�m���Og�H-�6fI`�RX0��RO�>4���-�;czk�
�K8w{H�
 �����9�hA���{�Kۮ�tw���k�Q�\>}�ҙ6L�e��:ج��n����,r�nt; 3���@�_���R����\�/�Y�mK�@
�V\��N.w�e�g9���JIz�c
�9�@��k�'��X��+����?qrM��X���"ǓQ�
9L��XLM�u_�T���5�����lo>sF�?�tf���i�:��fws�_�*�������v��Y;5�P{��i�d�H(��,Ǡ�bX� �A8�Lɘ냏��N�k|��W���ؙ�Yg�*��#��4�D"X~��y�:<ľ�uO'K>o��-�td���#-3��@wto�>�}�J��]$y�U�������,�d�%�¹���'�h�
yݽ���J�M��%�H�.���M�_�L�D�;(��'�s��j�qc��x��e	AGB�3q3�$�K���RMΖ��j�[9n�N�#��j���Pm�7��E�����YŧCE
��wH�����\HD{��#D�?ɢcq�;~���i�[It�	��|U5�$m*F�܎�`���E1�E��lC��?��)LI��!J&���l'�RK��N�����۶�!�������4��i�Y�6�L�o�����Ř���̭1r봽�t}Thm�t��^X�ʏ�1�d�<�N�u�H'F��J_r��D�i_�dќ�i��q�e�%k�Ƽ��"}�b�K�Y��8oȕ�M�r���0Yp��X��*=Ɓ����qmuSM=�e�\�R:�>�ӓbguv�p=�U�V�s�6��.V��Ar�s��Y��j��$!�j4T���
-��Յ�u�"1�i������s�Y���v�z�<����zA�y�6�9�p�nb�Qp�λH��]+U�h/���Rh��Q��zu���NCCg��}4 �n
���I���+���5"`b�WR3ҕ��F�o�L�W�5D��n�q_n�iw��)Wm�$�|i���4ϗj�^}�a��7Z�el�OM���h�=����b�0��g~�+N; c����.���]�\�h^h��r�dOF�33�&G{A�C������ ��e��0�����GX^i$�j���X�UL�I	ذj9�K��m�����}�=�M��'�ă��#b^���@\�AT�Ň!�}�P86�OPxv�4�^۔z��uY{�2�$o���3s֖2�O�����ӷ	2\k}�)�/O��j@�])�r�I�0�{���Zɲy����2�H\�܀3̘�����E4<�)��<9�Vo��Z��ǿ�Wg���#ŏ�ƮZ��I�Ǉ�i�H��ye��74�:WZ
��}O�b�Xn��ޒ�HK����*�m|X��A`�0[����9f�,l֒$X�V`,	�c�=S��0�8V�H�o���>̄�I�`��������9����ă᮷��G!C�4���K2��v�(z����na������쑧g�,�ƾ�q�ڠ{�tH�^�M3��7�0Д��e>`��[s)!�4�'�η�ד�x\�����|D�a2d�1RȺJcF���b���3�T��HS�0	�uQO��Ti&?�Ax��y���G1���/�fU2��c4`Ԋ��-ںVi�I2ZB>���6�ǜj����x,�d�ߡښL�TZw������}�wr��[!u�[=J��@-�h���k�n���b���:���d �p�N��G

'�丝�4E*c�?OYp�W7t)�s��ک,���&0��td��CU��)�՝k����^5^�;��R��{�W�u�߀��+7�M̹�A�Ǻ�l˘xu�r����<������dq6���*��/6�p�V��zSￔ=����g������@�vH���������T�{��� �����*L��A�E��?�K���Y�䋼Hu�c���ǒ��'�}ʔ==R�pku�v.�Q�WQN�"�O�4Cn7��Un��������m4�O=m�*
aB����=�P�߃L��"� +,ɴy�*��ñp*j><�%G��m�������r��L%N	ʶ�]R�*����D��#9��r	��R�:b�Ԓ��=�W�=d[�0L��ڏZ^��`�ݼ�շ`���ш��(""�yŃp[���
4
�%�3�m�f`�C
$/�j{昨),T�L�2Q�-�k7ԱS�EZs#�R�SvmE��X^�Z>3d M-H�ȿ��^��i�#��A<)v
�2W�V��q�3(衜BU�u�
b~0��!D����lv��Ȫ�]�
�q�6ww8ӺE���,[�kV���2p�y�V��H�"R$�#Ɉ��.a��%�^|�)��u%[�����: ޥ�f9���ÞJ�+,��x��saE����@���I��>�����P`���:�kg� N*��q�	k?� ��$���U5U�
�]K��0�G���e4v�ѩ��\fs��R��F�ɾ#�W)�.2m\G�D�x��V_1�󁮮V�6�ZRCXz�����ܝ�^_�-O��%�ke׌�N��l�{|�����zI�?�ԓ���������dr�[�vT��Z�Q�w^8~Q�\�:Y�t���]x���O`"M�k�	w��*cPa��<�
�����X��a[a�{8��{MP:�$s�B6�����	�v/�?�C�;�^��W�S�s�[�2���[\C��<xTl)��P60���.�"�-w#+����^	�l��p.�.'GBr��5�i�| ꩽ.d�E��,�ک��4<����xPpO��>P�7������)c��b$d�S��m��KJg/��.��/��v�k��uq�f�@y_��8تC��)e=��j�l5�e�T�2D�}yσa�\�;4�L����[nޜx�y�n�jÂ����Ė�H�.v���)��c@�9����#_[���7�r��e�YT'>��Ņ�qj1ܕ�Y����g�1g�^�sC7*�aMi��Q#�Bq@�J�
0�����,ƎF�2��Q���`��}X��w�Z�`Nw�^�fG�i\���l����/�t,��B<�0����E���oID�׼3��fs.V)Y�c_�]I�&q�����Oe�Z���<�9g�
 U��2���̙��I�½C���#L�K}�mVKt^����̓�K��EI��g��L�]L���-�aD���xg�����1��-t`U�0z]���xC�J�/1��v�����eп���ӵ3`�9fݹv.r��"Of@���� �9܂� @��)��B*�e�І��C�_����5��l�t�A����Pmmg�C����8�\5�ޫN]���Nf.�R3 ����	�^���Z�缥���t��������osE	M�"��]�D�B�Q��Iu��x^�N���=;��t�v;��1l��37�BN��xm����p�s������n��"����*T�A|����e�\��.��� U���:�[!��uD0{�J���iH���`q!J�T�9.��� 'R�F&0� w^m~�^�{�W�T�m���٣���*���{��O�X���z�1�� 
L�������C�G����/^��חX�(��� ��z���oAcRg� �zi��b��2-�Ry��$��m���Ȩg%���h�a��V��4#9;�gU�L��C��&	�`�Ҏz�*��B��>2Tɤ��xY�b�%3�ҷdn��8+޾`�s,���i|�4�.���/��B�	˂x�a�	�i)!H�{=>���w��"�
��߷ͪN#ϰ:���.����'a�µa�� p�<	��f3N�	��,�$RC߿&���� �?L���x!�Ex5�P���R� ¾w�+�/D���<>ϣ���a�+/8�'Y��h����&�*�b�k.�A�A�-��M�Q8��E��A]�FK91I�W"�ޫO�r�O���J�x��(�G�`k�L���Wk&��h~ܑ)���}��Ý,4
����J��4��.O��� ��3�YO/�+����{�0��++�ی���֍6���xTp�yĈF#�9�dD�C-!�/K���<j����B</	%;Z��m���<��"z��d�����+����俾3� ��2ḩ7��)zrG�d��t�oAK�c_�l>阶D�^?����0K���y��Fe�%9�.(�A`^��Fe�<�U���|�0�fM"�@,T4� @^/^��t=�mڸ��i�B5V`�|�?��Sm���U�OS����ә%�YS,.�� B�`.�Qs���2����`��bQåY�x�_,9���oc�%��e��u�Ek5\zs��f34)�UG\馒%�Ҟh��|"R��d9iD�+bT�{���;�HyQ]�9a	�l��%0fU����02g+��Y��Lg��D�bˣ~3j
"g��8]�	᧟e�xv�0
��
����ʭ"�gЃȰ���DI�%�3a��J�YUо=���T4йl2��͹������P��.L����{�.�����ݹ�RN���5���).#9���O�I\�'wϰ�����D���El�at������A��kܰ7�ֈh�+Ś�k4|cy��r�������Ow?ȸ'bCZ����kɣ�(El=٤޾"�ZUu�V�������6��U���GfUI�#R�38�5}�/�z��$������Wx�]��zn曏�ï>jx3[,����O%�4N$q��=��"���6��Ũ�}�����h�-L����H�M�����}�3�f���b>ݹ��ˊr�z�
�lA���]����N�\�V���"�lٜ�'+�$��_]f��&��^��<X����7qc��=�r�S3�bR�=�.�p���v���j0=dU�Q�Kp���}�}�L���k�f����o*��D�0��@IO͗˝�)e	r��	��]��m@�OYJ �K��U�e&�P�J�k[I�nTRЄL���k�g7�ځ)E]E�8y!���'�ae�
/=$���s�� �¤����L�lү��������C+��Lhc�_F͆s�����������z.j�C-M-�^��J4�����˞3�SZK1>5��¸�u4^*��ų�|���w	�73�(�n��?���2 �&6�Z��zTS�uB���ZҒ�������M5��ϒ34��̰��7�W�%�z)����t��m�l|!|֢�{y�L�וkcB�C����֓�u��= ���\��,�:��V�-c/_2-y��NBA�n��J�����)�v�Ty��]�Ih"�9��Jz&ë���������L�	Z�Y����lGs��`���y���r]V��+\K�NU�!���5Oͤ�g!A5ʡ*��\�5~�O[�H���AapŶ:͋m2���ZR]�y}�%�7sC:I	��%g�C�GL@>��"갖T9�B�n�)Q�)�2�M��M�� H�b�8XOD��2��p�`p3=
��tȝQϣB�����笠�҄�A&5��D
S{X�oG����Qٵ���� u)���kᲳN*�%��#Deh(�!=k�:��dIM<ݡ{\���6N�{ �IW49fW��Ƞ������]�G�&�rn���������)��+`3�G����nP>�7��9D%�ǌ�g/ ҅�UN�����-F*1� �,_�yoc�t�e���0�j�P��߷N)��7�8�]>d�˱���F�;�#`A{EH]tc��`I:x�p�o� *�&ޮϼ�7���.y�Nl)�1Ԏ=�n�'���b��o3F��r}���
��K����� {���,�)j���F�	匡o���a�L[��1�(�j�F�S,�7E�{�=��7?���D�z����� �!N+��eh�"L0���m9p�5L��.������Zt�һ6T�p�YE	�B�.H?���(Ѩ����?����v !��Ȧ'M�l�(ʋX���8�WQ�x�hʵCx���)������Yhe��(�ȝæZ7�a,f}!�"���~�ݎ�<9�H�38��E=�s��|O�R�ك���o� ��p��� �Gc�S�_�#��&�M��id�0�?
�\���WP/Ck��.zBT�����x�l=�c���B��Px�)�s�����X�ć�ұMƹ���®7�o�_��>�����o&��k��?B�8�z�h�����E��l�M�'B��֕�����`�Zp��-��|K��&�u�!�ϙ;��O�C�D��$&�kP��*�p0��E��&wQu���m��~W�W��w�,H�t�ÎY���0��L��+�	8�r$�y�9��R�K����������?�Q$$�gt�%S�;����Ù�論�jS椧�
�u�����*"t�����cf�Qn+�/�.��-���)`hdLm��9�,��Ѫ�4BW����`�' ��h�!��C�>�~��J@�`���t9���4l"�8UP[Ѕ��:��U�%�ŵsA�:�(�䇬���x�]��g8�+���oF_���R�A޶7�Y�3���R��R��Mu�x�o+�@i�j/�R+Lg+��`ՇS�L_����rLw^a^���W<��R#�?5�������M�na�6��w�v�~d�J]D�	JP��G�Q�
DZE��"�߾A�&��ve[5�OhE�K���ۛYy.��/N���DT��S����*�㐴#߸�yW���H��?�^�_�}�! �p�ug�e�`�.f&�hT'҉�,1�m<<]i> b���y�R����	��[U�f�P��i
��ܞ�C d�831#�OΩ!��ّ���n%Db���Z� �}��*���݃X1��4H�*�}�@FK�d�JR�@��& H�|�z�⇯�r_]���X�c��∻[��ԝ���>x���"�L=��F���^���U]�4|5BҰ���3�,Lx�pg�!Ss�2�Tq���P��1 �[B���Ѳ�z)�aIL�#	䯌�������i@h��(Z�?:���Jj z��:O.$��-�E���~@D$m<������˪���Qj��&f�6|��=�s���r�?ذ4bˇ�4����a]�[!�]a��r�唄�D�8,|�c�^N3�UYծP��):-�<�:��Kݍ}^�Ӄ1�}�a��Pt�T��j)a1zi�)2L��5����@�U��AYЋ�?��-.���7�>|oV��ղȭH0��h����<�m@��L�x��'M]^&��p$�]L�,���������)�}�P�g��»�35��R��Բ������2n�V:���;C� ��B���&ee�Az(Q�J�^�5(�؎�b�y+����Uv5d�zl3�z,wbBȪ���.�*x��wu��Ȏ��2?fBn��$?��/kG ߊr���_�z=�U11����"��C`>x�2y4��m���n�H���O����p`]��Q��si����*��RR�%G�Y'`�v����%��\�N�COg�86��z9�:ڴy��J����gwsW/��=��鬸��� E:t�a(�ͣb���v��"h��1$:NX��^���x/x�ϣ)u!uR9���?�$��3,��d�~�Y�k�/��V �2T�%f�wH���wCMw��EEnn��]"j��>�ħ��2�qO�R�vIYٌTiX�vÜ>��Q*$ ���H9���[�`�������o.��V/Ui��3Zx%�@T�AL���eW�� ����r"~��C�S��;�I��q[�n�,�$$C^ߖ��,F������.>]8�4�8�"�N��r�駿~��T6�tޝ]x�����Э��x��u�>x��,ٷ "���eH[���,� ���A�%���N|�?�[a�׍�u)*�Bڋ������tm�g�}G}G�� �p�`+��Sy�����Fc+:UܬW����W��������݀���sQ���1��¾-B5�d���l-׽����P�X��bbw�K�-r�kb��]]_�X<H?m�.��+N�F���i`�ŀ�M{����{_��Ͼ/*�l���G�/B�|��ݿ��M���� Z2���2��.�*�Ԧ�3h��K-�AБ&tf�gaޣhC��	�wp	js��Z�̱��5���1�pt�|�R�=�na�ҝc�c]�dZա¯"�b�mp;?�n$8jhn��!�-%Qm�����J�R�K��\��)���c�$��W��%���p�)�$�u��3L9W�Xy6�'p��v۔P?CKT6A;�E`cMD#O�GƇq��؄��b[�ʍ�kA��v�T�B��^4�S��?�d]8H�N_)1�j�s[kRL��7"��m�Bۀ=��o2d!@Ct}��6j��?T���(�R;|���/�����I�
��U���I;���d�~��-
���?��W̛dX�<�	��>�S��6b���2�M8�8P��'8�o~CfvY���X�|d|ܖ�ZT�m�z�-��f��'���oyZ#�Kq5��Y�/���x��j��q��H��@�wͥer�բ��eӤ���r�5��f����v��h��r��\�ۈ6�h�<�<�&�pq��aM*L����l5��I�T�s
�(���7t�v��O� ��5��2�Kx����e�q������7$�(I�x>Ò�h[MpP]��"f���i�����b�(� �kT�JC)q��kQdj͋G#K)�Q��>N8�}��1���s������s����7ʜ�[R+:`�`����w<+V�LdC����#&�铤-9hc���R�SR�5��d.�։>B/�B��Y��y�s�X�z�Վ��Ƀ��Mő�� ��qO)V3v�X��h�� ��^�	yJ�!N|����i�}0���ϲ��V�T�1خ)-̮�h�/����.Bĝq�|�+��l/����.�Zwv��\�$��?��:�,\h%�b��|S���~��7h���;f>�]��:�a������p��Ş�	Ud�Y���]�ar�,,P��Z�q�|/�� ]�z���eV�5*ˍ��±��)�&�;��ՏB����z�8fC�eĭ���V�#�l~��Zs��|��Q�.�1Le��g3�� ��dƸ�3�����Y?̦sv#��1��M�w
,�����X{���g7a\by9���$�V���,wݖF��d2qP2|���|��*��^6B�pL�ǫbig���+t�u�Dc4b9�����Jb���� �h@C��A8�VV�f?���z�2z�;F�,�����E_��-�g�M���MԲ�c5�(Nr��*�7q
 �%rQjK�5���e�M�H�d�'~J�U�oV��B��98iU�`�ڭ�Z�Y�f�L�TӜE�_d�ۻY���eUG�Z�x?�Q
��-�X���+���S@��Y�ȋ:̿����2�����~���HU�D�X����uj�:��,D\���gY"� �G;�YTnc	l��Iõ�Pљ�pYOr�q��m4���F����m����[L��E1$3Oaa<�$�%$f$|�t�Q/{؊D�2 �q�����6E!հ`�dG�{���dL'˺F-
�Ҝ]�	����� 4�.(Q[n9h"���KF��b�/���a��E�~��퀅�������3r�2�&o#쿫ߋ�������K�[~��h&��PЫ�(�Ҟ���<����x��dI�1�;;|��XI�m��).��_��@Y  :�X5�j���c5?��#҆�%yP�-�)t�U����+����0<<,���ӧz�EN�Tկ���a�n��KNi��v\�$�s,�fAN�R�͂��
�&n�}nHj���2�?
S��W }M�e,��8I�&Z�mGm�:��o��m"v�"�19K��V'�o��ii*I\Rc2���.�[&W�N���7P�*�En��Pmu��0���NVi��<��Q���v�	ҥ���8���?�Q�sw	d �i�J҅�UQ}qD�4-}B�ТA���`t�Ջ��x�:(Z<T<�(J� ��Y?|](���7'�y]O� �Gӱ�BhC��_ħ�o�{��"�e���L��*���W� V�q�sc�dT�;�\|{BT��W����z�f�����
��$����IgQ/��`17� }z�W�����p9A�!O�M�)ˇ���^f+�S�d�CR��){/ٴ�HNԤo�ױ��C���j���K"�D��U$�b����o���%�;��(��3��u�Ds�����,%�z:O�Z�KĶ@��gQr�M����NϠ�,�	s6�e9X ��������N���=�t��g��T���Ip���h��^�P�z&zc;~�Ue�3cY��y{?<Y�F�~��T��D��MŇ!/���>0V�iy��+Y�QٔA���z��C�[�C�eݼD�ZKz!��}������z���5o1��x�QXӻh�����C���d��'�(!M-Cм!C�5�QI9Dș��c�7=YՈ[,��m=o��k��aO�����]	�c���T=Y�ΚK)ʆ����6-s�e�~V�9�7�{k��5젇���)׈�S�zWQ8�w:S�ܱ]ގ�j �P��R�6�� ɧe�鸂&k�jOOeTl*��>�,3��*.�����*u�!�n��"�"c�;������ i��_$?k�\���Q%���v�x������et�Z�'���
ο�����](�2&᯵Y�'|Z���q���c�d�&�D���	#�fQu9a��D�$�_w��̽�'��S�`��f�[>�e��K���.f.���IY�����D�I/۽�H���'�pn�H�1p4(v������'��Y{�[cmjQE��5��s�UO�0;���ۨLM���s��~-;��j����7]��ꬣ[����r���Y��9;Ĉ	*I�*�'��7n�R�۲��G {��*�aF��D�0�	� ����)+$�قƤ�G��Wy�����M�ڧƶ�<U�7�B�z.H����"�ҟ��g��Gx�{@��P5��nĵ
����@��R�UAv6�������uS�}k��*�14-��`�3�^�Q�%��E"�V�s�c�R����́&�*av&�J�����Bн�
��Q��Y`�xE"|jb�J�/���B��v!�|���(���Tb�"�O@���ºw$t�~mR�a�ߘ�Isj{`��hE�ίL��p���?XC���Wxm?�uW�5E��B��ȸZ��!~Жs�;�^1��_��a�guQ�n�lx�1�99���.;���L4�TFLl�yO���-�o��p���t������AmNôPף�UMFJ{5�v��Rƌ;������@��@�@�^�q�|���P�aW�&N�e.��}�
$�E������e_=3�i�X2C,xQ�Z��)&B�1�[_7 utͅ=��3 �Br*��l�'���	b����S�l�d� f��8�N����$���ͯC���&Hy��'D�[������҄}b���� ��~Y�]��� ��/�f���J����ر�u�t�{?���8�?��ծ��J»�W.��k�&�[����aq�fs�J��̘\�Ԇ��;I.BZ/X-$�G,��a���U�!�W��i��n�д8[��8<����t��n��/q�؆�ٯԂPg��%��2�s�1L��_���^o�$\��a��h���L_�f�����m�qD>6Iq3V��8���@e;�&3,Yd�"L'JR��?I�fo������$��D�}}�[*��(�D�w��\��X� gc��`$j�>�W����W����T�"!_FC���4%n�b��X��9!�C{����Is,O���8g�]����b�ٞ�y�r�@~��NĒ�c�蒝�L�<�y��b�,�r�1�]�o H�H"> p]}�k�qK#z�;�>�B���p�#t����z
�lb�&P;3<4���I������6.%��sem��.�
��$ ��=t�x��i�?��}����˵p��B{6�{�Y;��(�Q|s7�[5��t��E��ߚ��J�k�FQv�e2�4���6ᛶ�ۉ�� �J���Z)8��\{���N�g�y�]F��e��"��i85�҃�AL7��/�t2�$�O�|6�����M��|�̱G��&41\u�4'�f�w?qf���M�F7r4m�-�wo@��j�Zʥ=���p=��ܛ ��@�%�+o��U���<�8hc�lͯlr��lҬ�N��Y�L�y�W��{�({Ѧ0���sd'=<�c�_��0~j݈���w��1��������F�Ղ�k&Ȩ1��5��z��Ԥ\PI�`_k�\�(�^o�ܡV�т2���$�����g:)�}%��oH���]�za�Q�g�n ���B� I����}�,iﯤ�y�uB�;��}�2�_!B��ɥ�h�"<ڋ]�a���u��D��ƺ`瘪*�ޘĸG�ڤ_v~3_KL��7z�� nm�a�#6�m�/�~B�!��U�˓��R�sbs��I�~�|�{����
|�&G>t�zd���GIU�5f��x�fd�Z�9�=±"��1�20�w���u�7x�\��"X�Q`b]Τ�Y��)a��P��_�ʹk���a�$F�/�� k�ik2D|{�3���@�Dr	�7|��O��\
j\e��b?g�jM��f�>~ڧb�*«��8tOb"�k�!�yQ�;<zU���l��/v0������I�V�q1�D���q�Ԟւ	%��B��v���x�"�c�o8K�Ϻ� u�߉B)�=�rF|�|JX���s�;�Gp$���!����?'��>�Ħ�&D�TA=���A?S/�� 9�1#?\�z�;R9�sG�-�H�����[�t>�loKÎ��^��'xXS	߅&L�V]����T��:6X?E��a�'��P��2��JU>7���=�mJŝ�d�'-�#h�
|�I�ށEc3�Z/�/d^�M�Ld����i"�}%�,��ވ�\!MvS2.��I���;$����.�3����H�y�w�����6�^��;��xg �1<�1�Ң��Z���*=�1v���Y�t��LK��Ss�E���k�@��@5�z\u���^�;%~RG���^�4P�p���I���A�2�R(�4�q;��h����1����M���6���:V���n�n]Tj���ËWթÊ�=o�!��mp.,0c�q��kG_�������W�X���a���83΄�m_�zF8Q�$��V������Q�	����C�%u��`�ٌF���Y��#�R<�jB?�n����7�j[��aT"�yh7rt��IfALE���k���]�^@��Em�!�²O�J�n��F����W�	�6���[��,v���j��A% ���l����a���keV'�����Z�ak�XH�o�r���:qiJ5��jJRhI��B���)�!J�0��<o��K(L�S�����@�[. 4�b͗��Qf�e^v�a��?0��,�RȄ����'c���*)e"5g?Q���@�ow��BJ��@�S�P���E�"�_D�����FD��>e�q�SiH�Ԃ)4 �)�L*'�+y��*��&gaXA�1l�-��a:3��{��ۆ2�N�$$q��}y��Zs{��$���2;p�p���S�Tkm���ڂp�����鄟
ǰ�N't�����������y��G[)�3�}N�9�~�Z}�Uv�?_�{�+��%l�֢D+��~�h�_�8i��io;��NP���rPc��;T�Ѯ�-	׹w�
�"nƋ��K�49����V+�JFc�^U�Qu�fq pt}
��"[h"��$�e�z�س=�)O�����9ӓVEi��zdd�5O��@�	2�ż(T��=��L�S!��u	�E��m�Ww�U�Z����n��g�Sa�|5��՚���G�������N�ny���D�e�sy�w��%t�]�UR+�	�&��A�$;9*���
%OM�o4b4����i�eA����`��N��=W�!���Io��v�*��b+<�:6��UH���N�\��ce���	�ryRd�eGe\CΫ�t�/X�K[+�#ϭ�|�W��R�ZԖ\����e�[�Ŕ)�J�>΁�fgo�k���1�b�}x�h$��&��:��:���DeXs�ǐ& Z�Hϣ+^��V/���}��'R�]�vп?�!Bo���:�R����#b�:Y"u�^�=q�M�e��Z�����Eך+�O����`@���CSѪE������hWP����8�b���Ď^�D�THim��B����hN\+�UP<+70"������h���g&�<�1��@����'����75������F�~�K/fW��`���#m"Wf��f��o�vr�NacU8���O$��\�{��{�(�|B��Mg���.q3"pj,��mⓋ|��/O{+(�@u]c�om7�ø��}�G_e�BP�>ʷ`�3c��ú%����VK�^Y����&�����@}�)V�7���>�fqP����� � �vK���5z�ET�'����.Ms&{Ş���d]��	�!���N"Ô��ۺۈ������X� �OXt���"�U�њ�� Ph�$��I�M�f��J[K��}A"4�5R�>�@���ޅXy�@
�y4���j���$P���4F%�eaF<��5�ő�]v��׵f�5� ��yV6�MF?��*l,�{:�K������G�Ǉ�]��k~��Sr��lAa�:���R��&p����;�U�:`��O�4�EjcPl��m3nI,R��׎>�5��N�N��o��q��T��	0�"�D޶�՘x$c�9�� ~��"O����&�T��i�A��o�[�q�$J�(>���eT䲝.���k�HT���3��u��g��aF����g�i8���6��=8
 ��s� 0)���
�6���9�+��=��{�I%�]P�RN!�����Ή0��!�yĜν^tK�6��^����Ȭ� YH�����I����7��Bw��%��I���E�޷�.��v�	zA3s{x!؆k���(�i����(p��M��1E|��a͟S��:��!��z���|�=�	�\�ʭ��LQ7 �T-Qw?�Z.ƽO?���n:;��U�!æ����FwȸN���5>��o˥m�0K���Y�Ft7o{���h������6�{�aH
��!1�zy���XH�+�0���V����r`�<��[�S������+�T��Fx�͏�L�@����R��>*�\���\�F~|.�D����)C�5���ib�i"m�Y�'�i��'��u,�7�GT��Ax�"P����"�_犡0�S-YO2�f��~�	�{#
3��#{S���ɪ�8C�s��}��3<9�Zxe�~����wg���e�RD������`�uҝ���	gv�7��ѧ!j�OC?��T�C6��d06`��LX$?�g�aȩ�S4���fM͘�p(����V-wS�_V!�0N��X�6�U�(h�z[܆��k��"����m<���h���^�,ͱL$��tv�� Z��+\�Edv�rz[��7���t��9����M^��E^��1r%'�:s3G��P�3��5grc�{h7W:�e��;�Ya=�QQ�:	��C�YF;J�_M8d�xj~�I�+f���𞷒�]V:�SH��g�[F8����M�v�����ucU���A>C؏I�&@�e8�x��)�-�ޒ���H��u ��7Pu��:����L$W����i�>�_x;�������p[r��� ���Y_i{+��p�Ʒ�����ĄX7O��+W,[������z�(�_2"�#�wN���/x�0&D	�8ϕ�N�jr$G���cp[1.9��E��K�H�eRs���ɣ���YL�7c3U|�k�2����L��q���4�J�hv��m��:�Y��ጥ�tP�/�B� d��#y�r1��e�R^2�j��>F�����M����y�#.�a�.d
�mf_{��p���m}`����)��}S7�C��g]f���N*�d���=����Q �z��>274ޙ�J0��#m�����W�Vz�o��!b�{�R��~�t���!��{Aj��:	AT5d��(��ꍍ&_�R)5R$݅�&�Ⱥ�+~�DY�z��]���/�=���F�߀ͤ��kC��=[�'uà@?i������_��c`Y��|��sT����ڐV�Y�՜Y�	�!�y4��P��;�Wp�HZz�ky}� ���9�YN�/9���_��zf>�:f�L^+S�4G�5;)[v)��r�������G�U��Т4��5k�Ӱ ��a�3�a�Vz�cuM�ck�K����X��9|�@/�ړ�9�hE�Dd����l�A?�l�O"�����l�@��c4V7�~�<�#�sUi��̿�`t�T% 5߰;s�F�әm-�R�M�0s0�!��.��s=��`E��i����X���E2|`���	�ׁf�~���gwDb�f�����uN���Z����=NeJ������\LJgX����Y8��|��!��u��~T���I-�T+�/��� ��_Ҍ�tS&���+��@�Q�o��째�����F�t^Aq�B�����]����9�S�p|����HąP�|2~{0���2�r�����ۺ�cF����vnyC�v��)ϴ�l�C���M�q�8ƺ��W��P�!3����^���)*�+�n��,�+�砜Dnu�׫l�軧C����>�eO�#�>%��_t�%\%	D�F����%7eπbI<��wb��vȺ���_ {M��B��9�l�|��g���S�� �;M���M�H��ܑ�;���Nf����Q@��@��x"yɤ^�,����t�9�h	(�"��d�KGa�]	� p��"�D�_�ny�Ȝ]�������Գ�H�$�\a;YA���L��CUT�L�,��d$t�zQ�#ѯ��=�O|S���k��4�����<P�{�q�$����j�������n�NY���]�Ū��sS�[�Ϲg�h��q��w��3�6{��ќ2; �a��-��}Z�_�%�N�<7��+�}�rC��hP��,o���>M����x�߬09J�0I���Ӻ���7O��T[gD��/���MG�E0���C�K S� fl.V;��,�v�Y	8�gr-`��C�G͒lY4Hl
�y�d~� �W�(!� >�*v˃1MT�I=�C&�)��f����r"P"Vb��	�gx��L�btR�b�gE�n��o~���%P�3�4�� ����]���z9���[��KCن��q�_#Qy`脗3<���]�H;0o�͗e �VIn'w�b�t\�R����D+O� �V��7|�K^$f�y��p �NZ���g!myz�i*��`�9ԁ�X�Yts��r�~����Y��x�n���͸��\S��^��WP���-��6����k<�|o�R�H�0�V7�.�&�:@�W����'MUeq������f��յt�EM`΍��-�(�G<z��(v�0�lߕ��$���+v�?dY����>��<��	y�1�����f��LO�`DEJ�_1AʐYD����R��ز�y��)�wjTq4=�%�V�s�5]�� �#��.^��ԑ�z���o���[S��]���\1ÅGx��؛9���UN�}���j�M3�y)E�.(���_�$�2̂_��̄--�4�^y��pϮ���q
B�u�z�;N�$,3,��as�������L���%t ���H.�%�%)����KT�g�oX�����)_3(���!�F��D���M� ��դǺ�`�@ǌ�	 ��ҭv�4� �8��ǋ�t����ǜ��Jq�\.�&�=��6+��1X;��ߦ���Fй��=����i�z�FP$�M�rS���L��i^����$s\R46�|�{�DUW�����{|�A�$x�~��!b�A���̽Z�r�~�x�����-|�,T���P����p��r��"�u���f�M��u��I��)�C�S!�E}	��j��>�������|wS=cX��X�p�)Y�I̒A���3 �I�F:�81�o���ʥ*n���}��"�l8u��I�y���n��Y���'�I��������*���7��' c���9�LVQ�I�d��T�;�'P�6_۽\/2�X9��|��5�p�}�Ka�����v'*U����9���j���3���WD�Ë2�\D_Hh7���Fyf�[�C�?�
�N"'�m3����0� >cu��u�y;�����_%� `U��6��[�#ޚq���G��k�̅���LF��0O%\@�c9G�����O]"�-�2�9^�FXN�ӊU_S��]UU���lD0�|��o	C����D�{	�sU�k�>��g)�+Y.���
8O�t�i��'G�QI"�����ے�\��Q�́C�A�4�`$��Lfj�.�vH[�͍�U"���]<�q�MD���n4�cI<@Ge��kPv�#��(~�$a�݁�A�'��.�U}�p�P�z�%?�T�&�I)�]*��g��^9,H��z���9o��(��/�܇�S�JNt��@XO<�
����2�]q�{v�$�d�H��U�<�\4��*�d5�m�L�5�P�臝H���ѥ!С#>R�s�cG�5�^~dh��=e��p�I�`s�d����19���h���9idr>?�B�*c/x2	ĵŐ�?&u���ł.�+*"�J{'� ���e��E�=��pM��K�{5�>N��U�m$�*s$S�D�x�E'KGK� �����K�8���������������C�]h�eqD7�G���ȷ�#m���d�����$�qݔAV|B��3��8(��H�LL���E_qJ���ˁ&��i�unw�[��.ס�a�F!eT�>�;�Jy�;�z*h� �kI�V�n�}r�����6����^Sc]�`:�s+���Id�_OͩJ-��˰Lr��+?�lpZ�/w�I���)ŋCMV�S��a�p��3�ST���>�瘉�������T`��P�@
l���(��۰��^_w�"o�}w:�ɿ����8،!�ȼRL3U�J���N�I��aг7��0�2�K�DŨzEк���zD�6-N��~#�P�����I/F�[�:Jh�B\�jđ|������V�{�z����kV��� ��a��!,�N��+^ �T��0���y��I��z��⹢�)GWaP�_qeb���FPWU��+_]��\�%1iL`��i�#�=����nE���V~��߳L`5�AìO��VEEM'v�F����$q�����lǓr�����h���}�����Ӳ,6"��sˁ��)wԘs`�4�A^���o���������n#t�}�ՁdеӧȊó�'�+��]����_��v�g��s����Kӕ�&�/�0s+]H�/��i����xme��,]�r��<����8�[\7<�'s.�k0�z���Ei{��������z����&�U�|�m��D�ǀ�ɟk��WA���u�q�9���F�=%�~��^8���4��f���������Y�����(���q�"�ܺ,�?P	��`�Z
T;Bڡէ�B������4|_ђ	/z`�˻��]�p��uR�l��f�p��'�����|�=�:ٜ���C�ӳ��N�1.W�\��9S"���B�8'���@�*<4��ͽV	���V^�vQyzŚҐ<��a	��X6�/���\�3�����8�ѷ���y�ʆ�W�5���+ض�� ���S.	�]�H.F^s����
��f!�MKR�1�ՠ���#E�}i���������3}Zi�2J?�S�sr�8��&�@�\������Is|f�#���o�0��,�ϡe�UGB��������Q�oX�kOT�G	w������N3���!9#���h17p�_k�}�x�k:gĽ��
\ |	�ߡ��E�G	puX3����.M/5�Nϝ~��!���I	��U-�@�)��5�okթ�
#qc���m�yg�RҠ#~�[��BO,O���]��%��2+�����}�<f��]p-�ڧy�z!���c�_>���Hͷ�J:Z�D��ikL�m����E��?�Z�z4A�B�|�מ����ɝ��t�jirQ���_���su½�t�=�2��(�$�ǆ�	�p=�����9�y�-2c��� W��;�@��"؆��0nV���5�&Ǒ:�.�.�J!]�7x$_^,��� ��dGZ���0z�:�/p5X�t�)��� �!��g6ݝ=� �
�d!md�����._g5,��򞃾\�'{_��޿Cy\�=��In�뗲���榱�@�o<>����	aV57�y8�2��|î��mq��U���:��}
@����`��̸-(�&��됪m9��v����j/�D���P�1��4'Q5c���]������W����pϣ5���A�Q�18b��W����g���� �l�N�|r��sÈ��B�p,�0�PV�A ���bF�eǌ�����
�_�+�3%��5^B�|�"�5Y�P�&��g�DWQ�]t*�t�Q�E�!Mi�n�J��gp�τ
ZC�G]��j�-�ښ����vtv�S�� S�2�zM&'L=��jJ&K=F&�-�>p���N;Hu��{��O��M�)E���SoKbx��pV�֜�*,����"�kt��z�1�WX�o��]f:G�$����u�L;�<=�~���,�U��Ӻ�����Fj,�
���HMD��c�,�:��W��X����l�h4k�]�8�M�����8R}ו@H���&�e2Ӑ���(�/h���C�~c9���tQ���#V ��t�!8�[FV�YڨX�J��|:�b���^�(�m�Q���'b.Q]�R���I���d����@�)ߙQ�u�u��%`�U1��meu�cR��4XZY�ஏ�|�ީA��Ħi�܅�I�؊��2j��U|m����$.@"-�����@�R15�"c��D4�T�Q���������b�/�L/ХH:�.Yo�%�7�B��z7P��ł45s���ו��G����1�D��h�xE;O��_�������87�0 5z���y�S�p��CLH3U-��N���;#�K�j��*�\ �$#�n����$Z���L�́��p�E����M�Z�{������z3 ���$A�����j"V�qxt�ąBQjaP�����$@�%cT����o������G"":��,X�	ax�7G�@���D{;z�B�ѷ/:$�L����_��ܰ����M!H��CuXk�vÍ��W>�5���b�h-/��zBcbS��,���4��t�B*:���Ŋ�Y��8E�c!���Z)���}�*tqMě���B�M�5�;�p�Vi��B�[���=��t<�z���d�X�t�g�ٗ�:��B���c'-d�Қq������tM$k�I��p����v�#rVW\F��/�}E�zV�N�����#�����z̈e#�a��i\~������RQ~�[�( Ʉ�L�?*꿛c|π-��z@��q�[i�rp���՜;���U;&v��P�='��Sౖ��|���sy$�����J+,a�y����%�o���C^���Hɒ[��FLct�|1!���=�����i��B>�`��ޗ�t��(Bg�1�a�Os�yh�Ӗ���۶�m��\��<�S�y1���@`$r��G{@��*s����7����x�}s
{�U�3;�X�X�A�!L�T+'��!�91��A輞e,Xg���'��}��y:u]�:�x"�8sr�^����9��v�I�4�o?F.����s��N�4L~�/ВTI�C��}'�,�<E5�)H��*�=��U�A�a�<:�9<W���\>ə�B��b
��ǷS���Wߴb��,�0> �����[�@m��N ���;�mH9Mףi�m~�nھ䷠���K��@G �J�D�&�V�d{���_��Z���x��H֓��q��W�)����汉����ӭM'��ޕ�U<��_O�5��QA��qY�tKJ�Έ�io݆�q��!�|cüF�Z$LkRG])����,�<N��}=/�_�s�I����o~���.�~)I>7�5�G5>F�ص�JF���7��l�K�h��Y+���T�']�1..Z�{�,�e~��+6��捎��Q�>v3-����C�]�s�2��R��e ��*½�����8^l��g�;�?e�25ӕ�TS8�pKzѧ�h�/)�D� ���~#�"���U�VȽ����O#�i.�R��W�k�q����osP�q�)�nHml�Ǖ��,/j���|a�r�����Zw����v����I�#�l+��S�����{|�-��R���J���|�Y\����)zT��/�<�?����R�	�Ž�
���HJ�3����~����AzP��N���0�Z���U���Jw4z-	�J�ӊFh�aR�ҥ�.]��K�T�\8~��z�� � ��m@��ț�y0�R u%:6�ӻ�O���3|��~�p�}��iKϵ��{)9�-��N�R�����}����Ë�.�)�j]b� n��ȇ"u�bZ�|�\��q��bBFH������i�,"�Tc��@pl����� �����ƍ?�Q6���D�=	����Sdy��a��N����4D�S����_���*��k0�%��&c,6tB�ӳG�/M��hL�2���j�%��C̅>���=� �t.�)Y�|&�ۦrK�W\�6��i��kv�[/�v�{܇��3�"�_Bqn��^�f��h��#�e�:�n=m�Ƚ�"m�j��Mɵ�VS�Yi�GX6��V���>�~+|�wJpKcY�\��nM��l�dF-�x_�Ì��:�:��_�P�傠�#�Q� m�x0���h�����5�!A�Y�b-s�`�P%��S0�(t���J�n~���>@�E%eU��Zì�`�� �Q_��KG+I7�4uB@���9Ո�H����.�
���e�:�-�>u�����n�4d�����QzO�P@��oqKתT}��/���0YJ�M��.em��(]T�Ս��x�&`k�Z���^6_TB���-6�*ӗ5n�~�������)�@������%�6��1'����[�U^�Ȥ}�(�->�b 	w�bm-� �ͲJ 5�7r�_dyR���j��8v��Ap��Ke��q/J�����{����ןq6��O?�������
W�= �kk�i��V<5j��|i�4�y����o��6X�8�r�t%�0B)��H0�K��;�z���ڣ��[��7�����f��Bӗ�yxCh�1�K=q
�*X5�k�&ً�i} � �.{�ɶ��I�ݸ<5���-�����#S�Y��k���}h�bAM8ڳ�a�~"y��<��m�A!+�f���hs7=B�R���lKj��b�Gn�jr��QS�FZ�{]�;����{���a�Y��"�"??�����27(�A�R����_ā�� nP��x]O˒ި䴓������?�z�.LO#${��d��(,gkE�b���J��&���9@�6g�<�>�JE�M�zo&�v~3�#A��c�\��k�
?�u�-��V��6.]���6&�[u�Yi�l��>ߍm��.�6Mߒ��!���jzϱ���#G���� �~�DK�B�.����q֓��b?.yඕ���Qt�r�����S/�ր��I��&��)���.�7�u���6�#���K�ԵZ5aH9��������� a��pr9az.�t���X��4o��h}����E(rgc^t���c���L��w�d�:.�� &�Ak�e�6l0¡@>���AT�5]*�b$����-V^_.Yq�9���
X���g�cf�v�@�Y6�����%g�`d�����nE��i۩!s�Ƹ>����k�O�6O��V�0�1v�Ð4�{`ΑE���:։d� ��cG2_�c�^�/�p�@����K�K�8w�sK)>���-"��v'�f�F��/���>/��S�9�����y�;��N8�;�cS�:�kEe�v2TȮ��O��"����O0q[�n'^�9s��e�؂Bk��X��6 ��K�� -G���Ɵ��c��Cq��-���G,E���P;M�2�D4q+g"'|Z�����9�u�=m�[�� ]@h1 /H�m�_���]��	dj���Ō�4����+vTR�s����;���v"�R[�5���a�T|r
�	>�0�J�ŝ4	'GP�y��0:Z����^+���ػ�\_�4g+���z`Y(�}S��ΝF+����(�r�w��'����<�G�� b�?�J:�����tP��}q�5\�C``#I<��ь݃���E^?G#a^K�D9���f^��o�%�6�$X�U*�2TP>	��R��T�`��%H����9��Oc�'�ȏA��1sj��e9��u�ڙ�	�yS�}� ���\�������'Gz�_j�#�G6��w�W8�uL�c[�c�s�����r֑�]}�l{sR�IPk.c�Dd��6mp�lW��^4�]��4�	���b��������'�K�.h�)�=����|�@(��?@�4�	o��0/%����{�-2�L'ˆ`�������$~#8�k".1g�!���2�FǞ�n�5G������X
�>q�68�^�=�D�)�v��'�aw�!���#ա��.!2أ�h��9�l~�X��9i�o�"��0�z�J�Zn	�/h��.�p{Tnd+.�qu�+���"��$�vc>.[k]%r�z��򋃹�]��)>��.��G�5��0ݱ��Z0�-Ԙt~��"�B�B���O�zL�A����u�d��v?e/�hp��K��JT]Zz�:�:�o{�"&����x���Z�u0.���d҄O0���_�#3��&�-^nI���� 3L���Q�����_�=�g�Z
�i���;��3G�:�l�Q9aW��b6���� ���+��WnP�(��p�V]�֥I�2��k�r��;b�����*I2��J�/�Ɵp�͑]��V�KX��H3��C�ޠ_ݹ�s�'�v�t���ᔈNob�^s-Y�h���s�z������:y�+��;����0D�(����&~1���"iρ(�Y������?�� OCW�S�YSe�������J�ůt��2��v�vƬ�֎�ƽ�����/̎f�t1܋�R�њ!)�lJC��Ov�@8r,9�b�0���eUB$s��8v�?�����";���0ʀ�|�F�����O���R��r�8��!�p;v�5�jy)�Z��{�Ż������{�~ps����υ��r�g7�ݠ!@�r��m#��=��'Xb( Mكz`JM���N'����p}��v�+�[MaG��=B!�u!mTq��xo8v�}̝m'����|�`�^J�l��g�+��� �Mg���G
�d�ׂ5����D�|��ޱf������}_��k�aC�l��h�n�<�\&��GR�_�<�6��,&�q	B���Y�ݾ�H��B(���p��v~�ĸF؄��/�Z/m���(��5������7"��0��E�ԏ،�0=�m]���1�v�#'�=X����r�Z���Q�����tԽ5F���i���@��6�&��;��]�\�߃h�Z@���R�Lݏ�e-�k5P?�6�yO�p+�����*�hU2CF��g'jo!鋃�TіRR�i,Z�T���S�����P��Eae���� 3�pK�#ZN��״���%A_��M���Y��"r} (��ɟ]mթj��D;��IL5'�ð����@�Ķ���9�xYc�
���-7^mw׈��y�!����
��#9��J�Ɇ����
������T�|<�Oakz�G~��������u��p��8(~L}��P�E��㎺a�Qonf��W���w�-8��`\�6P"=!�Y�̦]{/�ʀO�^�M��9e$��\d�YM�>!S�P,P����-�r��5eO�W�*��~%��틝��JB8�T١ˇ�(�<�`ɛ��*��)��$f��t���c����р䔴�#�]��?���6f|� a�C�bLN`_4�/��o�g~eA��ƚv�0�KV�LIF�����9xԍ�9��*oR�lO�Ey�A3�&���b~I}�)N��^��2����3���V��	7�����洖���b�N>��ӭ���.܉C땵^�avS�d�ZS�Ouw��Gª��+�H�W�Q�����ãFỈB���T]C�7Q�1@���+h�o95T�W�@�pC��3�	������'��p$躋$����"|���j�t��;]�T���AnvFD��f$��u���u�"�UА�1�����W�o����,�p�c���{Yu%�o�Kҏ>٢gA�n��JG��V�̥M�1֋j�p��R�᭔�O<��!q^TEp��k��(�х�8�������MH&R�����1�+�%_�huw�l��>�(��Ň�i�v4�X��Z�}�����[4j�"���!_(���ˬ��-�[�1��twHG�p�6~L־��-j��{����!q;x������/D��mB[&�nb��3pDY!�n�8\*5�Ĭ�c��+
��_�4:mȐ��S9�FX-�� �r�#��1��n��l�� ���:�e�C���&z׽k��=1g)���y��[[ua����7�EH�R���,��/&J��ު���B����#�+I�r�҄���B����\P���)B�I��Wt!��qg�o�}����{ZHo��w!�;i
�w�hs����ȹ~�b���&#��e5R"X[��w_�^���|������dX6�+z.��d4g�
[��F�ّ�8��~7&��
���4��^�N���_��1�E�G�����$À{KT����X��I$�HBrUO�qE��5��P�K.��B,��N��5�����M�vj]�[���-�	��z�e+T��#��M4�q�!��9b꥚P�W�����ho�����^0��L��'�cI�0�`zē�-z�� F�I��	�v���g�q�3]��)��o_�ɤ �*t��%�O�I�\G�æ!'�f�է4<+�`:�,��Ze�%
�����	]��G2&ج�����ȼ�'�Bz��
��}Ŏ�˻A���9sނ�5^���UO~����1c��5�=E.��GV����v@o����x䧱���"����h�#F�y�\�$D��[<7~r�sM��E�u�����%��<���%�~�1E�1VZxV�TK?U���.e0Y-ϓ�sO��8{��	�3��Dh�-j�Z,\��N�m�Ux�}4�3�G�@����5�G���)k�F��L1%�ķn�q^�Ը�N&�uЁ�$����:�@y�*-��x�]<�+��iL�W���P��֧�.�H5�7f�'ILeM�pon4w�AD)���er>��O�Y���
�*����hf���Z#v�%z0�
:[
�=�QO�Ølp�r&�� `U� ���3�|�%R�:P�F�
� �W�Slt�R�$i6����\h�Y���!�L��mQ��q�Tĭ�Mr����h����cO#�$�'�cNI̡mL�J�
����Rn|���zI���:����. S���s�瀆���|C޲L��k,��h���rl!Da�����(��J:�lk�ςv�v�u��	������!H��ŕM/&@z���_x��Z����d`����D������@J�a�ʄ�,[	p��e^��,��`iʷ:�<���YY���Y�s� �t��r�4{~$�by��ҽ��*t�tF3|�B>����m�Io�����M�<]��_zPa~5�f2<�ݟ�epD�z�p��A�B��a�!��9�s���½<覂����Ϊ$0��N���~�Ma��s�ogEK����]�BC΄�븪��n�6"��3��@��=C�(�&	�L��lө� �]��=�g]�l��,�˞C.�J���WWv�w ��]ϷD���x9.��9(��Wc5���k6�MN"��te��i��[�ꕡ���%�Q|�	��4{�j�j,��a�;���t#Q�r,3�}"����Ԯ�dM� ��D��]�D���,�����H���$�lS��?)1�(����e�:�Ah�M&��v�}=��&�!���4֑���C�v�z��Hs3�|�l��c'4��3��|p��vC�擌���&��f�H�(V��_E�J�R&,�&�H�?ƹ{�=��V/?���VY-<I�==��i��з) ۼ��9�	��(�_���U�O{)��`e�E��g�q`3�